/*
* Copyright 2019 International Business Machines
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*/
`timescale 1ns/1ps

module gqeJoin_wrapper (
    stall_start_ext,
    stall_done_ext,
    stall_start_str,
    stall_done_str,
    stall_start_int,
    stall_done_int,
    s_axi_control_AWADDR,
    s_axi_control_AWVALID,
    s_axi_control_AWREADY,
    s_axi_control_WDATA,
    s_axi_control_WSTRB,
    s_axi_control_WVALID,
    s_axi_control_WREADY,
    s_axi_control_BRESP,
    s_axi_control_BVALID,
    s_axi_control_BREADY,
    s_axi_control_ARADDR,
    s_axi_control_ARVALID,
    s_axi_control_ARREADY,
    s_axi_control_RDATA,
    s_axi_control_RRESP,
    s_axi_control_RVALID,
    s_axi_control_RREADY,
    ap_clk,
    ap_rst_n,
    event_done,
    interrupt,
    event_start,
    m_axi_gmem0_0_AWADDR,
    m_axi_gmem0_0_AWLEN,
    m_axi_gmem0_0_AWSIZE,
    m_axi_gmem0_0_AWBURST,
    m_axi_gmem0_0_AWLOCK,
    m_axi_gmem0_0_AWREGION,
    m_axi_gmem0_0_AWCACHE,
    m_axi_gmem0_0_AWPROT,
    m_axi_gmem0_0_AWQOS,
    m_axi_gmem0_0_AWVALID,
    m_axi_gmem0_0_AWREADY,
    m_axi_gmem0_0_WDATA,
    m_axi_gmem0_0_WSTRB,
    m_axi_gmem0_0_WLAST,
    m_axi_gmem0_0_WVALID,
    m_axi_gmem0_0_WREADY,
    m_axi_gmem0_0_BRESP,
    m_axi_gmem0_0_BVALID,
    m_axi_gmem0_0_BREADY,
    m_axi_gmem0_0_ARADDR,
    m_axi_gmem0_0_ARLEN,
    m_axi_gmem0_0_ARSIZE,
    m_axi_gmem0_0_ARBURST,
    m_axi_gmem0_0_ARLOCK,
    m_axi_gmem0_0_ARREGION,
    m_axi_gmem0_0_ARCACHE,
    m_axi_gmem0_0_ARPROT,
    m_axi_gmem0_0_ARQOS,
    m_axi_gmem0_0_ARVALID,
    m_axi_gmem0_0_ARREADY,
    m_axi_gmem0_0_RDATA,
    m_axi_gmem0_0_RRESP,
    m_axi_gmem0_0_RLAST,
    m_axi_gmem0_0_RVALID,
    m_axi_gmem0_0_RREADY,
    m_axi_gmem0_1_AWADDR,
    m_axi_gmem0_1_AWLEN,
    m_axi_gmem0_1_AWSIZE,
    m_axi_gmem0_1_AWBURST,
    m_axi_gmem0_1_AWLOCK,
    m_axi_gmem0_1_AWREGION,
    m_axi_gmem0_1_AWCACHE,
    m_axi_gmem0_1_AWPROT,
    m_axi_gmem0_1_AWQOS,
    m_axi_gmem0_1_AWVALID,
    m_axi_gmem0_1_AWREADY,
    m_axi_gmem0_1_WDATA,
    m_axi_gmem0_1_WSTRB,
    m_axi_gmem0_1_WLAST,
    m_axi_gmem0_1_WVALID,
    m_axi_gmem0_1_WREADY,
    m_axi_gmem0_1_BRESP,
    m_axi_gmem0_1_BVALID,
    m_axi_gmem0_1_BREADY,
    m_axi_gmem0_1_ARADDR,
    m_axi_gmem0_1_ARLEN,
    m_axi_gmem0_1_ARSIZE,
    m_axi_gmem0_1_ARBURST,
    m_axi_gmem0_1_ARLOCK,
    m_axi_gmem0_1_ARREGION,
    m_axi_gmem0_1_ARCACHE,
    m_axi_gmem0_1_ARPROT,
    m_axi_gmem0_1_ARQOS,
    m_axi_gmem0_1_ARVALID,
    m_axi_gmem0_1_ARREADY,
    m_axi_gmem0_1_RDATA,
    m_axi_gmem0_1_RRESP,
    m_axi_gmem0_1_RLAST,
    m_axi_gmem0_1_RVALID,
    m_axi_gmem0_1_RREADY,
    m_axi_gmem0_2_AWADDR,
    m_axi_gmem0_2_AWLEN,
    m_axi_gmem0_2_AWSIZE,
    m_axi_gmem0_2_AWBURST,
    m_axi_gmem0_2_AWLOCK,
    m_axi_gmem0_2_AWREGION,
    m_axi_gmem0_2_AWCACHE,
    m_axi_gmem0_2_AWPROT,
    m_axi_gmem0_2_AWQOS,
    m_axi_gmem0_2_AWVALID,
    m_axi_gmem0_2_AWREADY,
    m_axi_gmem0_2_WDATA,
    m_axi_gmem0_2_WSTRB,
    m_axi_gmem0_2_WLAST,
    m_axi_gmem0_2_WVALID,
    m_axi_gmem0_2_WREADY,
    m_axi_gmem0_2_BRESP,
    m_axi_gmem0_2_BVALID,
    m_axi_gmem0_2_BREADY,
    m_axi_gmem0_2_ARADDR,
    m_axi_gmem0_2_ARLEN,
    m_axi_gmem0_2_ARSIZE,
    m_axi_gmem0_2_ARBURST,
    m_axi_gmem0_2_ARLOCK,
    m_axi_gmem0_2_ARREGION,
    m_axi_gmem0_2_ARCACHE,
    m_axi_gmem0_2_ARPROT,
    m_axi_gmem0_2_ARQOS,
    m_axi_gmem0_2_ARVALID,
    m_axi_gmem0_2_ARREADY,
    m_axi_gmem0_2_RDATA,
    m_axi_gmem0_2_RRESP,
    m_axi_gmem0_2_RLAST,
    m_axi_gmem0_2_RVALID,
    m_axi_gmem0_2_RREADY,
    m_axi_gmem0_3_AWADDR,
    m_axi_gmem0_3_AWLEN,
    m_axi_gmem0_3_AWSIZE,
    m_axi_gmem0_3_AWBURST,
    m_axi_gmem0_3_AWLOCK,
    m_axi_gmem0_3_AWREGION,
    m_axi_gmem0_3_AWCACHE,
    m_axi_gmem0_3_AWPROT,
    m_axi_gmem0_3_AWQOS,
    m_axi_gmem0_3_AWVALID,
    m_axi_gmem0_3_AWREADY,
    m_axi_gmem0_3_WDATA,
    m_axi_gmem0_3_WSTRB,
    m_axi_gmem0_3_WLAST,
    m_axi_gmem0_3_WVALID,
    m_axi_gmem0_3_WREADY,
    m_axi_gmem0_3_BRESP,
    m_axi_gmem0_3_BVALID,
    m_axi_gmem0_3_BREADY,
    m_axi_gmem0_3_ARADDR,
    m_axi_gmem0_3_ARLEN,
    m_axi_gmem0_3_ARSIZE,
    m_axi_gmem0_3_ARBURST,
    m_axi_gmem0_3_ARLOCK,
    m_axi_gmem0_3_ARREGION,
    m_axi_gmem0_3_ARCACHE,
    m_axi_gmem0_3_ARPROT,
    m_axi_gmem0_3_ARQOS,
    m_axi_gmem0_3_ARVALID,
    m_axi_gmem0_3_ARREADY,
    m_axi_gmem0_3_RDATA,
    m_axi_gmem0_3_RRESP,
    m_axi_gmem0_3_RLAST,
    m_axi_gmem0_3_RVALID,
    m_axi_gmem0_3_RREADY,
    m_axi_gmem1_0_AWADDR,
    m_axi_gmem1_0_AWLEN,
    m_axi_gmem1_0_AWSIZE,
    m_axi_gmem1_0_AWBURST,
    m_axi_gmem1_0_AWLOCK,
    m_axi_gmem1_0_AWREGION,
    m_axi_gmem1_0_AWCACHE,
    m_axi_gmem1_0_AWPROT,
    m_axi_gmem1_0_AWQOS,
    m_axi_gmem1_0_AWVALID,
    m_axi_gmem1_0_AWREADY,
    m_axi_gmem1_0_WDATA,
    m_axi_gmem1_0_WSTRB,
    m_axi_gmem1_0_WLAST,
    m_axi_gmem1_0_WVALID,
    m_axi_gmem1_0_WREADY,
    m_axi_gmem1_0_BRESP,
    m_axi_gmem1_0_BVALID,
    m_axi_gmem1_0_BREADY,
    m_axi_gmem1_0_ARADDR,
    m_axi_gmem1_0_ARLEN,
    m_axi_gmem1_0_ARSIZE,
    m_axi_gmem1_0_ARBURST,
    m_axi_gmem1_0_ARLOCK,
    m_axi_gmem1_0_ARREGION,
    m_axi_gmem1_0_ARCACHE,
    m_axi_gmem1_0_ARPROT,
    m_axi_gmem1_0_ARQOS,
    m_axi_gmem1_0_ARVALID,
    m_axi_gmem1_0_ARREADY,
    m_axi_gmem1_0_RDATA,
    m_axi_gmem1_0_RRESP,
    m_axi_gmem1_0_RLAST,
    m_axi_gmem1_0_RVALID,
    m_axi_gmem1_0_RREADY,
    m_axi_gmem1_1_AWADDR,
    m_axi_gmem1_1_AWLEN,
    m_axi_gmem1_1_AWSIZE,
    m_axi_gmem1_1_AWBURST,
    m_axi_gmem1_1_AWLOCK,
    m_axi_gmem1_1_AWREGION,
    m_axi_gmem1_1_AWCACHE,
    m_axi_gmem1_1_AWPROT,
    m_axi_gmem1_1_AWQOS,
    m_axi_gmem1_1_AWVALID,
    m_axi_gmem1_1_AWREADY,
    m_axi_gmem1_1_WDATA,
    m_axi_gmem1_1_WSTRB,
    m_axi_gmem1_1_WLAST,
    m_axi_gmem1_1_WVALID,
    m_axi_gmem1_1_WREADY,
    m_axi_gmem1_1_BRESP,
    m_axi_gmem1_1_BVALID,
    m_axi_gmem1_1_BREADY,
    m_axi_gmem1_1_ARADDR,
    m_axi_gmem1_1_ARLEN,
    m_axi_gmem1_1_ARSIZE,
    m_axi_gmem1_1_ARBURST,
    m_axi_gmem1_1_ARLOCK,
    m_axi_gmem1_1_ARREGION,
    m_axi_gmem1_1_ARCACHE,
    m_axi_gmem1_1_ARPROT,
    m_axi_gmem1_1_ARQOS,
    m_axi_gmem1_1_ARVALID,
    m_axi_gmem1_1_ARREADY,
    m_axi_gmem1_1_RDATA,
    m_axi_gmem1_1_RRESP,
    m_axi_gmem1_1_RLAST,
    m_axi_gmem1_1_RVALID,
    m_axi_gmem1_1_RREADY,
    m_axi_gmem1_2_AWADDR,
    m_axi_gmem1_2_AWLEN,
    m_axi_gmem1_2_AWSIZE,
    m_axi_gmem1_2_AWBURST,
    m_axi_gmem1_2_AWLOCK,
    m_axi_gmem1_2_AWREGION,
    m_axi_gmem1_2_AWCACHE,
    m_axi_gmem1_2_AWPROT,
    m_axi_gmem1_2_AWQOS,
    m_axi_gmem1_2_AWVALID,
    m_axi_gmem1_2_AWREADY,
    m_axi_gmem1_2_WDATA,
    m_axi_gmem1_2_WSTRB,
    m_axi_gmem1_2_WLAST,
    m_axi_gmem1_2_WVALID,
    m_axi_gmem1_2_WREADY,
    m_axi_gmem1_2_BRESP,
    m_axi_gmem1_2_BVALID,
    m_axi_gmem1_2_BREADY,
    m_axi_gmem1_2_ARADDR,
    m_axi_gmem1_2_ARLEN,
    m_axi_gmem1_2_ARSIZE,
    m_axi_gmem1_2_ARBURST,
    m_axi_gmem1_2_ARLOCK,
    m_axi_gmem1_2_ARREGION,
    m_axi_gmem1_2_ARCACHE,
    m_axi_gmem1_2_ARPROT,
    m_axi_gmem1_2_ARQOS,
    m_axi_gmem1_2_ARVALID,
    m_axi_gmem1_2_ARREADY,
    m_axi_gmem1_2_RDATA,
    m_axi_gmem1_2_RRESP,
    m_axi_gmem1_2_RLAST,
    m_axi_gmem1_2_RVALID,
    m_axi_gmem1_2_RREADY,
    m_axi_gmem1_3_AWADDR,
    m_axi_gmem1_3_AWLEN,
    m_axi_gmem1_3_AWSIZE,
    m_axi_gmem1_3_AWBURST,
    m_axi_gmem1_3_AWLOCK,
    m_axi_gmem1_3_AWREGION,
    m_axi_gmem1_3_AWCACHE,
    m_axi_gmem1_3_AWPROT,
    m_axi_gmem1_3_AWQOS,
    m_axi_gmem1_3_AWVALID,
    m_axi_gmem1_3_AWREADY,
    m_axi_gmem1_3_WDATA,
    m_axi_gmem1_3_WSTRB,
    m_axi_gmem1_3_WLAST,
    m_axi_gmem1_3_WVALID,
    m_axi_gmem1_3_WREADY,
    m_axi_gmem1_3_BRESP,
    m_axi_gmem1_3_BVALID,
    m_axi_gmem1_3_BREADY,
    m_axi_gmem1_3_ARADDR,
    m_axi_gmem1_3_ARLEN,
    m_axi_gmem1_3_ARSIZE,
    m_axi_gmem1_3_ARBURST,
    m_axi_gmem1_3_ARLOCK,
    m_axi_gmem1_3_ARREGION,
    m_axi_gmem1_3_ARCACHE,
    m_axi_gmem1_3_ARPROT,
    m_axi_gmem1_3_ARQOS,
    m_axi_gmem1_3_ARVALID,
    m_axi_gmem1_3_ARREADY,
    m_axi_gmem1_3_RDATA,
    m_axi_gmem1_3_RRESP,
    m_axi_gmem1_3_RLAST,
    m_axi_gmem1_3_RVALID,
    m_axi_gmem1_3_RREADY,
    m_axi_gmem1_4_AWADDR,
    m_axi_gmem1_4_AWLEN,
    m_axi_gmem1_4_AWSIZE,
    m_axi_gmem1_4_AWBURST,
    m_axi_gmem1_4_AWLOCK,
    m_axi_gmem1_4_AWREGION,
    m_axi_gmem1_4_AWCACHE,
    m_axi_gmem1_4_AWPROT,
    m_axi_gmem1_4_AWQOS,
    m_axi_gmem1_4_AWVALID,
    m_axi_gmem1_4_AWREADY,
    m_axi_gmem1_4_WDATA,
    m_axi_gmem1_4_WSTRB,
    m_axi_gmem1_4_WLAST,
    m_axi_gmem1_4_WVALID,
    m_axi_gmem1_4_WREADY,
    m_axi_gmem1_4_BRESP,
    m_axi_gmem1_4_BVALID,
    m_axi_gmem1_4_BREADY,
    m_axi_gmem1_4_ARADDR,
    m_axi_gmem1_4_ARLEN,
    m_axi_gmem1_4_ARSIZE,
    m_axi_gmem1_4_ARBURST,
    m_axi_gmem1_4_ARLOCK,
    m_axi_gmem1_4_ARREGION,
    m_axi_gmem1_4_ARCACHE,
    m_axi_gmem1_4_ARPROT,
    m_axi_gmem1_4_ARQOS,
    m_axi_gmem1_4_ARVALID,
    m_axi_gmem1_4_ARREADY,
    m_axi_gmem1_4_RDATA,
    m_axi_gmem1_4_RRESP,
    m_axi_gmem1_4_RLAST,
    m_axi_gmem1_4_RVALID,
    m_axi_gmem1_4_RREADY,
    m_axi_gmem1_5_AWADDR,
    m_axi_gmem1_5_AWLEN,
    m_axi_gmem1_5_AWSIZE,
    m_axi_gmem1_5_AWBURST,
    m_axi_gmem1_5_AWLOCK,
    m_axi_gmem1_5_AWREGION,
    m_axi_gmem1_5_AWCACHE,
    m_axi_gmem1_5_AWPROT,
    m_axi_gmem1_5_AWQOS,
    m_axi_gmem1_5_AWVALID,
    m_axi_gmem1_5_AWREADY,
    m_axi_gmem1_5_WDATA,
    m_axi_gmem1_5_WSTRB,
    m_axi_gmem1_5_WLAST,
    m_axi_gmem1_5_WVALID,
    m_axi_gmem1_5_WREADY,
    m_axi_gmem1_5_BRESP,
    m_axi_gmem1_5_BVALID,
    m_axi_gmem1_5_BREADY,
    m_axi_gmem1_5_ARADDR,
    m_axi_gmem1_5_ARLEN,
    m_axi_gmem1_5_ARSIZE,
    m_axi_gmem1_5_ARBURST,
    m_axi_gmem1_5_ARLOCK,
    m_axi_gmem1_5_ARREGION,
    m_axi_gmem1_5_ARCACHE,
    m_axi_gmem1_5_ARPROT,
    m_axi_gmem1_5_ARQOS,
    m_axi_gmem1_5_ARVALID,
    m_axi_gmem1_5_ARREADY,
    m_axi_gmem1_5_RDATA,
    m_axi_gmem1_5_RRESP,
    m_axi_gmem1_5_RLAST,
    m_axi_gmem1_5_RVALID,
    m_axi_gmem1_5_RREADY,
    m_axi_gmem1_6_AWADDR,
    m_axi_gmem1_6_AWLEN,
    m_axi_gmem1_6_AWSIZE,
    m_axi_gmem1_6_AWBURST,
    m_axi_gmem1_6_AWLOCK,
    m_axi_gmem1_6_AWREGION,
    m_axi_gmem1_6_AWCACHE,
    m_axi_gmem1_6_AWPROT,
    m_axi_gmem1_6_AWQOS,
    m_axi_gmem1_6_AWVALID,
    m_axi_gmem1_6_AWREADY,
    m_axi_gmem1_6_WDATA,
    m_axi_gmem1_6_WSTRB,
    m_axi_gmem1_6_WLAST,
    m_axi_gmem1_6_WVALID,
    m_axi_gmem1_6_WREADY,
    m_axi_gmem1_6_BRESP,
    m_axi_gmem1_6_BVALID,
    m_axi_gmem1_6_BREADY,
    m_axi_gmem1_6_ARADDR,
    m_axi_gmem1_6_ARLEN,
    m_axi_gmem1_6_ARSIZE,
    m_axi_gmem1_6_ARBURST,
    m_axi_gmem1_6_ARLOCK,
    m_axi_gmem1_6_ARREGION,
    m_axi_gmem1_6_ARCACHE,
    m_axi_gmem1_6_ARPROT,
    m_axi_gmem1_6_ARQOS,
    m_axi_gmem1_6_ARVALID,
    m_axi_gmem1_6_ARREADY,
    m_axi_gmem1_6_RDATA,
    m_axi_gmem1_6_RRESP,
    m_axi_gmem1_6_RLAST,
    m_axi_gmem1_6_RVALID,
    m_axi_gmem1_6_RREADY,
    m_axi_gmem1_7_AWADDR,
    m_axi_gmem1_7_AWLEN,
    m_axi_gmem1_7_AWSIZE,
    m_axi_gmem1_7_AWBURST,
    m_axi_gmem1_7_AWLOCK,
    m_axi_gmem1_7_AWREGION,
    m_axi_gmem1_7_AWCACHE,
    m_axi_gmem1_7_AWPROT,
    m_axi_gmem1_7_AWQOS,
    m_axi_gmem1_7_AWVALID,
    m_axi_gmem1_7_AWREADY,
    m_axi_gmem1_7_WDATA,
    m_axi_gmem1_7_WSTRB,
    m_axi_gmem1_7_WLAST,
    m_axi_gmem1_7_WVALID,
    m_axi_gmem1_7_WREADY,
    m_axi_gmem1_7_BRESP,
    m_axi_gmem1_7_BVALID,
    m_axi_gmem1_7_BREADY,
    m_axi_gmem1_7_ARADDR,
    m_axi_gmem1_7_ARLEN,
    m_axi_gmem1_7_ARSIZE,
    m_axi_gmem1_7_ARBURST,
    m_axi_gmem1_7_ARLOCK,
    m_axi_gmem1_7_ARREGION,
    m_axi_gmem1_7_ARCACHE,
    m_axi_gmem1_7_ARPROT,
    m_axi_gmem1_7_ARQOS,
    m_axi_gmem1_7_ARVALID,
    m_axi_gmem1_7_ARREADY,
    m_axi_gmem1_7_RDATA,
    m_axi_gmem1_7_RRESP,
    m_axi_gmem1_7_RLAST,
    m_axi_gmem1_7_RVALID,
    m_axi_gmem1_7_RREADY,
    m_axi_gmem2_0_AWADDR,
    m_axi_gmem2_0_AWLEN,
    m_axi_gmem2_0_AWSIZE,
    m_axi_gmem2_0_AWBURST,
    m_axi_gmem2_0_AWLOCK,
    m_axi_gmem2_0_AWREGION,
    m_axi_gmem2_0_AWCACHE,
    m_axi_gmem2_0_AWPROT,
    m_axi_gmem2_0_AWQOS,
    m_axi_gmem2_0_AWVALID,
    m_axi_gmem2_0_AWREADY,
    m_axi_gmem2_0_WDATA,
    m_axi_gmem2_0_WSTRB,
    m_axi_gmem2_0_WLAST,
    m_axi_gmem2_0_WVALID,
    m_axi_gmem2_0_WREADY,
    m_axi_gmem2_0_BRESP,
    m_axi_gmem2_0_BVALID,
    m_axi_gmem2_0_BREADY,
    m_axi_gmem2_0_ARADDR,
    m_axi_gmem2_0_ARLEN,
    m_axi_gmem2_0_ARSIZE,
    m_axi_gmem2_0_ARBURST,
    m_axi_gmem2_0_ARLOCK,
    m_axi_gmem2_0_ARREGION,
    m_axi_gmem2_0_ARCACHE,
    m_axi_gmem2_0_ARPROT,
    m_axi_gmem2_0_ARQOS,
    m_axi_gmem2_0_ARVALID,
    m_axi_gmem2_0_ARREADY,
    m_axi_gmem2_0_RDATA,
    m_axi_gmem2_0_RRESP,
    m_axi_gmem2_0_RLAST,
    m_axi_gmem2_0_RVALID,
    m_axi_gmem2_0_RREADY,
    m_axi_gmem2_1_AWADDR,
    m_axi_gmem2_1_AWLEN,
    m_axi_gmem2_1_AWSIZE,
    m_axi_gmem2_1_AWBURST,
    m_axi_gmem2_1_AWLOCK,
    m_axi_gmem2_1_AWREGION,
    m_axi_gmem2_1_AWCACHE,
    m_axi_gmem2_1_AWPROT,
    m_axi_gmem2_1_AWQOS,
    m_axi_gmem2_1_AWVALID,
    m_axi_gmem2_1_AWREADY,
    m_axi_gmem2_1_WDATA,
    m_axi_gmem2_1_WSTRB,
    m_axi_gmem2_1_WLAST,
    m_axi_gmem2_1_WVALID,
    m_axi_gmem2_1_WREADY,
    m_axi_gmem2_1_BRESP,
    m_axi_gmem2_1_BVALID,
    m_axi_gmem2_1_BREADY,
    m_axi_gmem2_1_ARADDR,
    m_axi_gmem2_1_ARLEN,
    m_axi_gmem2_1_ARSIZE,
    m_axi_gmem2_1_ARBURST,
    m_axi_gmem2_1_ARLOCK,
    m_axi_gmem2_1_ARREGION,
    m_axi_gmem2_1_ARCACHE,
    m_axi_gmem2_1_ARPROT,
    m_axi_gmem2_1_ARQOS,
    m_axi_gmem2_1_ARVALID,
    m_axi_gmem2_1_ARREADY,
    m_axi_gmem2_1_RDATA,
    m_axi_gmem2_1_RRESP,
    m_axi_gmem2_1_RLAST,
    m_axi_gmem2_1_RVALID,
    m_axi_gmem2_1_RREADY,
    m_axi_gmem2_2_AWADDR,
    m_axi_gmem2_2_AWLEN,
    m_axi_gmem2_2_AWSIZE,
    m_axi_gmem2_2_AWBURST,
    m_axi_gmem2_2_AWLOCK,
    m_axi_gmem2_2_AWREGION,
    m_axi_gmem2_2_AWCACHE,
    m_axi_gmem2_2_AWPROT,
    m_axi_gmem2_2_AWQOS,
    m_axi_gmem2_2_AWVALID,
    m_axi_gmem2_2_AWREADY,
    m_axi_gmem2_2_WDATA,
    m_axi_gmem2_2_WSTRB,
    m_axi_gmem2_2_WLAST,
    m_axi_gmem2_2_WVALID,
    m_axi_gmem2_2_WREADY,
    m_axi_gmem2_2_BRESP,
    m_axi_gmem2_2_BVALID,
    m_axi_gmem2_2_BREADY,
    m_axi_gmem2_2_ARADDR,
    m_axi_gmem2_2_ARLEN,
    m_axi_gmem2_2_ARSIZE,
    m_axi_gmem2_2_ARBURST,
    m_axi_gmem2_2_ARLOCK,
    m_axi_gmem2_2_ARREGION,
    m_axi_gmem2_2_ARCACHE,
    m_axi_gmem2_2_ARPROT,
    m_axi_gmem2_2_ARQOS,
    m_axi_gmem2_2_ARVALID,
    m_axi_gmem2_2_ARREADY,
    m_axi_gmem2_2_RDATA,
    m_axi_gmem2_2_RRESP,
    m_axi_gmem2_2_RLAST,
    m_axi_gmem2_2_RVALID,
    m_axi_gmem2_2_RREADY,
    m_axi_gmem2_3_AWADDR,
    m_axi_gmem2_3_AWLEN,
    m_axi_gmem2_3_AWSIZE,
    m_axi_gmem2_3_AWBURST,
    m_axi_gmem2_3_AWLOCK,
    m_axi_gmem2_3_AWREGION,
    m_axi_gmem2_3_AWCACHE,
    m_axi_gmem2_3_AWPROT,
    m_axi_gmem2_3_AWQOS,
    m_axi_gmem2_3_AWVALID,
    m_axi_gmem2_3_AWREADY,
    m_axi_gmem2_3_WDATA,
    m_axi_gmem2_3_WSTRB,
    m_axi_gmem2_3_WLAST,
    m_axi_gmem2_3_WVALID,
    m_axi_gmem2_3_WREADY,
    m_axi_gmem2_3_BRESP,
    m_axi_gmem2_3_BVALID,
    m_axi_gmem2_3_BREADY,
    m_axi_gmem2_3_ARADDR,
    m_axi_gmem2_3_ARLEN,
    m_axi_gmem2_3_ARSIZE,
    m_axi_gmem2_3_ARBURST,
    m_axi_gmem2_3_ARLOCK,
    m_axi_gmem2_3_ARREGION,
    m_axi_gmem2_3_ARCACHE,
    m_axi_gmem2_3_ARPROT,
    m_axi_gmem2_3_ARQOS,
    m_axi_gmem2_3_ARVALID,
    m_axi_gmem2_3_ARREADY,
    m_axi_gmem2_3_RDATA,
    m_axi_gmem2_3_RRESP,
    m_axi_gmem2_3_RLAST,
    m_axi_gmem2_3_RVALID,
    m_axi_gmem2_3_RREADY,
    m_axi_gmem2_4_AWADDR,
    m_axi_gmem2_4_AWLEN,
    m_axi_gmem2_4_AWSIZE,
    m_axi_gmem2_4_AWBURST,
    m_axi_gmem2_4_AWLOCK,
    m_axi_gmem2_4_AWREGION,
    m_axi_gmem2_4_AWCACHE,
    m_axi_gmem2_4_AWPROT,
    m_axi_gmem2_4_AWQOS,
    m_axi_gmem2_4_AWVALID,
    m_axi_gmem2_4_AWREADY,
    m_axi_gmem2_4_WDATA,
    m_axi_gmem2_4_WSTRB,
    m_axi_gmem2_4_WLAST,
    m_axi_gmem2_4_WVALID,
    m_axi_gmem2_4_WREADY,
    m_axi_gmem2_4_BRESP,
    m_axi_gmem2_4_BVALID,
    m_axi_gmem2_4_BREADY,
    m_axi_gmem2_4_ARADDR,
    m_axi_gmem2_4_ARLEN,
    m_axi_gmem2_4_ARSIZE,
    m_axi_gmem2_4_ARBURST,
    m_axi_gmem2_4_ARLOCK,
    m_axi_gmem2_4_ARREGION,
    m_axi_gmem2_4_ARCACHE,
    m_axi_gmem2_4_ARPROT,
    m_axi_gmem2_4_ARQOS,
    m_axi_gmem2_4_ARVALID,
    m_axi_gmem2_4_ARREADY,
    m_axi_gmem2_4_RDATA,
    m_axi_gmem2_4_RRESP,
    m_axi_gmem2_4_RLAST,
    m_axi_gmem2_4_RVALID,
    m_axi_gmem2_4_RREADY,
    m_axi_gmem2_5_AWADDR,
    m_axi_gmem2_5_AWLEN,
    m_axi_gmem2_5_AWSIZE,
    m_axi_gmem2_5_AWBURST,
    m_axi_gmem2_5_AWLOCK,
    m_axi_gmem2_5_AWREGION,
    m_axi_gmem2_5_AWCACHE,
    m_axi_gmem2_5_AWPROT,
    m_axi_gmem2_5_AWQOS,
    m_axi_gmem2_5_AWVALID,
    m_axi_gmem2_5_AWREADY,
    m_axi_gmem2_5_WDATA,
    m_axi_gmem2_5_WSTRB,
    m_axi_gmem2_5_WLAST,
    m_axi_gmem2_5_WVALID,
    m_axi_gmem2_5_WREADY,
    m_axi_gmem2_5_BRESP,
    m_axi_gmem2_5_BVALID,
    m_axi_gmem2_5_BREADY,
    m_axi_gmem2_5_ARADDR,
    m_axi_gmem2_5_ARLEN,
    m_axi_gmem2_5_ARSIZE,
    m_axi_gmem2_5_ARBURST,
    m_axi_gmem2_5_ARLOCK,
    m_axi_gmem2_5_ARREGION,
    m_axi_gmem2_5_ARCACHE,
    m_axi_gmem2_5_ARPROT,
    m_axi_gmem2_5_ARQOS,
    m_axi_gmem2_5_ARVALID,
    m_axi_gmem2_5_ARREADY,
    m_axi_gmem2_5_RDATA,
    m_axi_gmem2_5_RRESP,
    m_axi_gmem2_5_RLAST,
    m_axi_gmem2_5_RVALID,
    m_axi_gmem2_5_RREADY,
    m_axi_gmem2_6_AWADDR,
    m_axi_gmem2_6_AWLEN,
    m_axi_gmem2_6_AWSIZE,
    m_axi_gmem2_6_AWBURST,
    m_axi_gmem2_6_AWLOCK,
    m_axi_gmem2_6_AWREGION,
    m_axi_gmem2_6_AWCACHE,
    m_axi_gmem2_6_AWPROT,
    m_axi_gmem2_6_AWQOS,
    m_axi_gmem2_6_AWVALID,
    m_axi_gmem2_6_AWREADY,
    m_axi_gmem2_6_WDATA,
    m_axi_gmem2_6_WSTRB,
    m_axi_gmem2_6_WLAST,
    m_axi_gmem2_6_WVALID,
    m_axi_gmem2_6_WREADY,
    m_axi_gmem2_6_BRESP,
    m_axi_gmem2_6_BVALID,
    m_axi_gmem2_6_BREADY,
    m_axi_gmem2_6_ARADDR,
    m_axi_gmem2_6_ARLEN,
    m_axi_gmem2_6_ARSIZE,
    m_axi_gmem2_6_ARBURST,
    m_axi_gmem2_6_ARLOCK,
    m_axi_gmem2_6_ARREGION,
    m_axi_gmem2_6_ARCACHE,
    m_axi_gmem2_6_ARPROT,
    m_axi_gmem2_6_ARQOS,
    m_axi_gmem2_6_ARVALID,
    m_axi_gmem2_6_ARREADY,
    m_axi_gmem2_6_RDATA,
    m_axi_gmem2_6_RRESP,
    m_axi_gmem2_6_RLAST,
    m_axi_gmem2_6_RVALID,
    m_axi_gmem2_6_RREADY,
    m_axi_gmem2_7_AWADDR,
    m_axi_gmem2_7_AWLEN,
    m_axi_gmem2_7_AWSIZE,
    m_axi_gmem2_7_AWBURST,
    m_axi_gmem2_7_AWLOCK,
    m_axi_gmem2_7_AWREGION,
    m_axi_gmem2_7_AWCACHE,
    m_axi_gmem2_7_AWPROT,
    m_axi_gmem2_7_AWQOS,
    m_axi_gmem2_7_AWVALID,
    m_axi_gmem2_7_AWREADY,
    m_axi_gmem2_7_WDATA,
    m_axi_gmem2_7_WSTRB,
    m_axi_gmem2_7_WLAST,
    m_axi_gmem2_7_WVALID,
    m_axi_gmem2_7_WREADY,
    m_axi_gmem2_7_BRESP,
    m_axi_gmem2_7_BVALID,
    m_axi_gmem2_7_BREADY,
    m_axi_gmem2_7_ARADDR,
    m_axi_gmem2_7_ARLEN,
    m_axi_gmem2_7_ARSIZE,
    m_axi_gmem2_7_ARBURST,
    m_axi_gmem2_7_ARLOCK,
    m_axi_gmem2_7_ARREGION,
    m_axi_gmem2_7_ARCACHE,
    m_axi_gmem2_7_ARPROT,
    m_axi_gmem2_7_ARQOS,
    m_axi_gmem2_7_ARVALID,
    m_axi_gmem2_7_ARREADY,
    m_axi_gmem2_7_RDATA,
    m_axi_gmem2_7_RRESP,
    m_axi_gmem2_7_RLAST,
    m_axi_gmem2_7_RVALID,
    m_axi_gmem2_7_RREADY
    );

    output wire stall_start_ext;
    output wire stall_done_ext;
    output wire stall_start_str;
    output wire stall_done_str;
    output wire stall_start_int;
    output wire stall_done_int;
    input wire [7 : 0] s_axi_control_AWADDR;
    input wire s_axi_control_AWVALID;
    output wire s_axi_control_AWREADY;
    input wire [31 : 0] s_axi_control_WDATA;
    input wire [3 : 0] s_axi_control_WSTRB;
    input wire s_axi_control_WVALID;
    output wire s_axi_control_WREADY;
    output wire [1 : 0] s_axi_control_BRESP;
    output wire s_axi_control_BVALID;
    input wire s_axi_control_BREADY;
    input wire [7 : 0] s_axi_control_ARADDR;
    input wire s_axi_control_ARVALID;
    output wire s_axi_control_ARREADY;
    output wire [31 : 0] s_axi_control_RDATA;
    output wire [1 : 0] s_axi_control_RRESP;
    output wire s_axi_control_RVALID;
    input wire s_axi_control_RREADY;
    input wire ap_clk;
    input wire ap_rst_n;
    output wire event_done;
    output wire interrupt;
    output wire event_start;
    output wire [63 : 0] m_axi_gmem0_0_AWADDR;
    output wire [7 : 0] m_axi_gmem0_0_AWLEN;
    output wire [2 : 0] m_axi_gmem0_0_AWSIZE;
    output wire [1 : 0] m_axi_gmem0_0_AWBURST;
    output wire [1 : 0] m_axi_gmem0_0_AWLOCK;
    output wire [3 : 0] m_axi_gmem0_0_AWREGION;
    output wire [3 : 0] m_axi_gmem0_0_AWCACHE;
    output wire [2 : 0] m_axi_gmem0_0_AWPROT;
    output wire [3 : 0] m_axi_gmem0_0_AWQOS;
    output wire m_axi_gmem0_0_AWVALID;
    input wire m_axi_gmem0_0_AWREADY;
    output wire [511 : 0] m_axi_gmem0_0_WDATA;
    output wire [63 : 0] m_axi_gmem0_0_WSTRB;
    output wire m_axi_gmem0_0_WLAST;
    output wire m_axi_gmem0_0_WVALID;
    input wire m_axi_gmem0_0_WREADY;
    input wire [1 : 0] m_axi_gmem0_0_BRESP;
    input wire m_axi_gmem0_0_BVALID;
    output wire m_axi_gmem0_0_BREADY;
    output wire [63 : 0] m_axi_gmem0_0_ARADDR;
    output wire [7 : 0] m_axi_gmem0_0_ARLEN;
    output wire [2 : 0] m_axi_gmem0_0_ARSIZE;
    output wire [1 : 0] m_axi_gmem0_0_ARBURST;
    output wire [1 : 0] m_axi_gmem0_0_ARLOCK;
    output wire [3 : 0] m_axi_gmem0_0_ARREGION;
    output wire [3 : 0] m_axi_gmem0_0_ARCACHE;
    output wire [2 : 0] m_axi_gmem0_0_ARPROT;
    output wire [3 : 0] m_axi_gmem0_0_ARQOS;
    output wire m_axi_gmem0_0_ARVALID;
    input wire m_axi_gmem0_0_ARREADY;
    input wire [511 : 0] m_axi_gmem0_0_RDATA;
    input wire [1 : 0] m_axi_gmem0_0_RRESP;
    input wire m_axi_gmem0_0_RLAST;
    input wire m_axi_gmem0_0_RVALID;
    output wire m_axi_gmem0_0_RREADY;
    output wire [63 : 0] m_axi_gmem0_1_AWADDR;
    output wire [7 : 0] m_axi_gmem0_1_AWLEN;
    output wire [2 : 0] m_axi_gmem0_1_AWSIZE;
    output wire [1 : 0] m_axi_gmem0_1_AWBURST;
    output wire [1 : 0] m_axi_gmem0_1_AWLOCK;
    output wire [3 : 0] m_axi_gmem0_1_AWREGION;
    output wire [3 : 0] m_axi_gmem0_1_AWCACHE;
    output wire [2 : 0] m_axi_gmem0_1_AWPROT;
    output wire [3 : 0] m_axi_gmem0_1_AWQOS;
    output wire m_axi_gmem0_1_AWVALID;
    input wire m_axi_gmem0_1_AWREADY;
    output wire [511 : 0] m_axi_gmem0_1_WDATA;
    output wire [63 : 0] m_axi_gmem0_1_WSTRB;
    output wire m_axi_gmem0_1_WLAST;
    output wire m_axi_gmem0_1_WVALID;
    input wire m_axi_gmem0_1_WREADY;
    input wire [1 : 0] m_axi_gmem0_1_BRESP;
    input wire m_axi_gmem0_1_BVALID;
    output wire m_axi_gmem0_1_BREADY;
    output wire [63 : 0] m_axi_gmem0_1_ARADDR;
    output wire [7 : 0] m_axi_gmem0_1_ARLEN;
    output wire [2 : 0] m_axi_gmem0_1_ARSIZE;
    output wire [1 : 0] m_axi_gmem0_1_ARBURST;
    output wire [1 : 0] m_axi_gmem0_1_ARLOCK;
    output wire [3 : 0] m_axi_gmem0_1_ARREGION;
    output wire [3 : 0] m_axi_gmem0_1_ARCACHE;
    output wire [2 : 0] m_axi_gmem0_1_ARPROT;
    output wire [3 : 0] m_axi_gmem0_1_ARQOS;
    output wire m_axi_gmem0_1_ARVALID;
    input wire m_axi_gmem0_1_ARREADY;
    input wire [511 : 0] m_axi_gmem0_1_RDATA;
    input wire [1 : 0] m_axi_gmem0_1_RRESP;
    input wire m_axi_gmem0_1_RLAST;
    input wire m_axi_gmem0_1_RVALID;
    output wire m_axi_gmem0_1_RREADY;
    output wire [63 : 0] m_axi_gmem0_2_AWADDR;
    output wire [7 : 0] m_axi_gmem0_2_AWLEN;
    output wire [2 : 0] m_axi_gmem0_2_AWSIZE;
    output wire [1 : 0] m_axi_gmem0_2_AWBURST;
    output wire [1 : 0] m_axi_gmem0_2_AWLOCK;
    output wire [3 : 0] m_axi_gmem0_2_AWREGION;
    output wire [3 : 0] m_axi_gmem0_2_AWCACHE;
    output wire [2 : 0] m_axi_gmem0_2_AWPROT;
    output wire [3 : 0] m_axi_gmem0_2_AWQOS;
    output wire m_axi_gmem0_2_AWVALID;
    input wire m_axi_gmem0_2_AWREADY;
    output wire [511 : 0] m_axi_gmem0_2_WDATA;
    output wire [63 : 0] m_axi_gmem0_2_WSTRB;
    output wire m_axi_gmem0_2_WLAST;
    output wire m_axi_gmem0_2_WVALID;
    input wire m_axi_gmem0_2_WREADY;
    input wire [1 : 0] m_axi_gmem0_2_BRESP;
    input wire m_axi_gmem0_2_BVALID;
    output wire m_axi_gmem0_2_BREADY;
    output wire [63 : 0] m_axi_gmem0_2_ARADDR;
    output wire [7 : 0] m_axi_gmem0_2_ARLEN;
    output wire [2 : 0] m_axi_gmem0_2_ARSIZE;
    output wire [1 : 0] m_axi_gmem0_2_ARBURST;
    output wire [1 : 0] m_axi_gmem0_2_ARLOCK;
    output wire [3 : 0] m_axi_gmem0_2_ARREGION;
    output wire [3 : 0] m_axi_gmem0_2_ARCACHE;
    output wire [2 : 0] m_axi_gmem0_2_ARPROT;
    output wire [3 : 0] m_axi_gmem0_2_ARQOS;
    output wire m_axi_gmem0_2_ARVALID;
    input wire m_axi_gmem0_2_ARREADY;
    input wire [511 : 0] m_axi_gmem0_2_RDATA;
    input wire [1 : 0] m_axi_gmem0_2_RRESP;
    input wire m_axi_gmem0_2_RLAST;
    input wire m_axi_gmem0_2_RVALID;
    output wire m_axi_gmem0_2_RREADY;
    output wire [63 : 0] m_axi_gmem0_3_AWADDR;
    output wire [7 : 0] m_axi_gmem0_3_AWLEN;
    output wire [2 : 0] m_axi_gmem0_3_AWSIZE;
    output wire [1 : 0] m_axi_gmem0_3_AWBURST;
    output wire [1 : 0] m_axi_gmem0_3_AWLOCK;
    output wire [3 : 0] m_axi_gmem0_3_AWREGION;
    output wire [3 : 0] m_axi_gmem0_3_AWCACHE;
    output wire [2 : 0] m_axi_gmem0_3_AWPROT;
    output wire [3 : 0] m_axi_gmem0_3_AWQOS;
    output wire m_axi_gmem0_3_AWVALID;
    input wire m_axi_gmem0_3_AWREADY;
    output wire [511 : 0] m_axi_gmem0_3_WDATA;
    output wire [63 : 0] m_axi_gmem0_3_WSTRB;
    output wire m_axi_gmem0_3_WLAST;
    output wire m_axi_gmem0_3_WVALID;
    input wire m_axi_gmem0_3_WREADY;
    input wire [1 : 0] m_axi_gmem0_3_BRESP;
    input wire m_axi_gmem0_3_BVALID;
    output wire m_axi_gmem0_3_BREADY;
    output wire [63 : 0] m_axi_gmem0_3_ARADDR;
    output wire [7 : 0] m_axi_gmem0_3_ARLEN;
    output wire [2 : 0] m_axi_gmem0_3_ARSIZE;
    output wire [1 : 0] m_axi_gmem0_3_ARBURST;
    output wire [1 : 0] m_axi_gmem0_3_ARLOCK;
    output wire [3 : 0] m_axi_gmem0_3_ARREGION;
    output wire [3 : 0] m_axi_gmem0_3_ARCACHE;
    output wire [2 : 0] m_axi_gmem0_3_ARPROT;
    output wire [3 : 0] m_axi_gmem0_3_ARQOS;
    output wire m_axi_gmem0_3_ARVALID;
    input wire m_axi_gmem0_3_ARREADY;
    input wire [511 : 0] m_axi_gmem0_3_RDATA;
    input wire [1 : 0] m_axi_gmem0_3_RRESP;
    input wire m_axi_gmem0_3_RLAST;
    input wire m_axi_gmem0_3_RVALID;
    output wire m_axi_gmem0_3_RREADY;
    output wire [63 : 0] m_axi_gmem1_0_AWADDR;
    output wire [7 : 0] m_axi_gmem1_0_AWLEN;
    output wire [2 : 0] m_axi_gmem1_0_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_0_AWBURST;
    output wire [1 : 0] m_axi_gmem1_0_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_0_AWREGION;
    output wire [3 : 0] m_axi_gmem1_0_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_0_AWPROT;
    output wire [3 : 0] m_axi_gmem1_0_AWQOS;
    output wire m_axi_gmem1_0_AWVALID;
    input wire m_axi_gmem1_0_AWREADY;
    output wire [63 : 0] m_axi_gmem1_0_WDATA;
    output wire [7 : 0] m_axi_gmem1_0_WSTRB;
    output wire m_axi_gmem1_0_WLAST;
    output wire m_axi_gmem1_0_WVALID;
    input wire m_axi_gmem1_0_WREADY;
    input wire [1 : 0] m_axi_gmem1_0_BRESP;
    input wire m_axi_gmem1_0_BVALID;
    output wire m_axi_gmem1_0_BREADY;
    output wire [63 : 0] m_axi_gmem1_0_ARADDR;
    output wire [7 : 0] m_axi_gmem1_0_ARLEN;
    output wire [2 : 0] m_axi_gmem1_0_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_0_ARBURST;
    output wire [1 : 0] m_axi_gmem1_0_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_0_ARREGION;
    output wire [3 : 0] m_axi_gmem1_0_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_0_ARPROT;
    output wire [3 : 0] m_axi_gmem1_0_ARQOS;
    output wire m_axi_gmem1_0_ARVALID;
    input wire m_axi_gmem1_0_ARREADY;
    input wire [63 : 0] m_axi_gmem1_0_RDATA;
    input wire [1 : 0] m_axi_gmem1_0_RRESP;
    input wire m_axi_gmem1_0_RLAST;
    input wire m_axi_gmem1_0_RVALID;
    output wire m_axi_gmem1_0_RREADY;
    output wire [63 : 0] m_axi_gmem1_1_AWADDR;
    output wire [7 : 0] m_axi_gmem1_1_AWLEN;
    output wire [2 : 0] m_axi_gmem1_1_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_1_AWBURST;
    output wire [1 : 0] m_axi_gmem1_1_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_1_AWREGION;
    output wire [3 : 0] m_axi_gmem1_1_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_1_AWPROT;
    output wire [3 : 0] m_axi_gmem1_1_AWQOS;
    output wire m_axi_gmem1_1_AWVALID;
    input wire m_axi_gmem1_1_AWREADY;
    output wire [63 : 0] m_axi_gmem1_1_WDATA;
    output wire [7 : 0] m_axi_gmem1_1_WSTRB;
    output wire m_axi_gmem1_1_WLAST;
    output wire m_axi_gmem1_1_WVALID;
    input wire m_axi_gmem1_1_WREADY;
    input wire [1 : 0] m_axi_gmem1_1_BRESP;
    input wire m_axi_gmem1_1_BVALID;
    output wire m_axi_gmem1_1_BREADY;
    output wire [63 : 0] m_axi_gmem1_1_ARADDR;
    output wire [7 : 0] m_axi_gmem1_1_ARLEN;
    output wire [2 : 0] m_axi_gmem1_1_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_1_ARBURST;
    output wire [1 : 0] m_axi_gmem1_1_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_1_ARREGION;
    output wire [3 : 0] m_axi_gmem1_1_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_1_ARPROT;
    output wire [3 : 0] m_axi_gmem1_1_ARQOS;
    output wire m_axi_gmem1_1_ARVALID;
    input wire m_axi_gmem1_1_ARREADY;
    input wire [63 : 0] m_axi_gmem1_1_RDATA;
    input wire [1 : 0] m_axi_gmem1_1_RRESP;
    input wire m_axi_gmem1_1_RLAST;
    input wire m_axi_gmem1_1_RVALID;
    output wire m_axi_gmem1_1_RREADY;
    output wire [63 : 0] m_axi_gmem1_2_AWADDR;
    output wire [7 : 0] m_axi_gmem1_2_AWLEN;
    output wire [2 : 0] m_axi_gmem1_2_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_2_AWBURST;
    output wire [1 : 0] m_axi_gmem1_2_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_2_AWREGION;
    output wire [3 : 0] m_axi_gmem1_2_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_2_AWPROT;
    output wire [3 : 0] m_axi_gmem1_2_AWQOS;
    output wire m_axi_gmem1_2_AWVALID;
    input wire m_axi_gmem1_2_AWREADY;
    output wire [63 : 0] m_axi_gmem1_2_WDATA;
    output wire [7 : 0] m_axi_gmem1_2_WSTRB;
    output wire m_axi_gmem1_2_WLAST;
    output wire m_axi_gmem1_2_WVALID;
    input wire m_axi_gmem1_2_WREADY;
    input wire [1 : 0] m_axi_gmem1_2_BRESP;
    input wire m_axi_gmem1_2_BVALID;
    output wire m_axi_gmem1_2_BREADY;
    output wire [63 : 0] m_axi_gmem1_2_ARADDR;
    output wire [7 : 0] m_axi_gmem1_2_ARLEN;
    output wire [2 : 0] m_axi_gmem1_2_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_2_ARBURST;
    output wire [1 : 0] m_axi_gmem1_2_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_2_ARREGION;
    output wire [3 : 0] m_axi_gmem1_2_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_2_ARPROT;
    output wire [3 : 0] m_axi_gmem1_2_ARQOS;
    output wire m_axi_gmem1_2_ARVALID;
    input wire m_axi_gmem1_2_ARREADY;
    input wire [63 : 0] m_axi_gmem1_2_RDATA;
    input wire [1 : 0] m_axi_gmem1_2_RRESP;
    input wire m_axi_gmem1_2_RLAST;
    input wire m_axi_gmem1_2_RVALID;
    output wire m_axi_gmem1_2_RREADY;
    output wire [63 : 0] m_axi_gmem1_3_AWADDR;
    output wire [7 : 0] m_axi_gmem1_3_AWLEN;
    output wire [2 : 0] m_axi_gmem1_3_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_3_AWBURST;
    output wire [1 : 0] m_axi_gmem1_3_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_3_AWREGION;
    output wire [3 : 0] m_axi_gmem1_3_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_3_AWPROT;
    output wire [3 : 0] m_axi_gmem1_3_AWQOS;
    output wire m_axi_gmem1_3_AWVALID;
    input wire m_axi_gmem1_3_AWREADY;
    output wire [63 : 0] m_axi_gmem1_3_WDATA;
    output wire [7 : 0] m_axi_gmem1_3_WSTRB;
    output wire m_axi_gmem1_3_WLAST;
    output wire m_axi_gmem1_3_WVALID;
    input wire m_axi_gmem1_3_WREADY;
    input wire [1 : 0] m_axi_gmem1_3_BRESP;
    input wire m_axi_gmem1_3_BVALID;
    output wire m_axi_gmem1_3_BREADY;
    output wire [63 : 0] m_axi_gmem1_3_ARADDR;
    output wire [7 : 0] m_axi_gmem1_3_ARLEN;
    output wire [2 : 0] m_axi_gmem1_3_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_3_ARBURST;
    output wire [1 : 0] m_axi_gmem1_3_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_3_ARREGION;
    output wire [3 : 0] m_axi_gmem1_3_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_3_ARPROT;
    output wire [3 : 0] m_axi_gmem1_3_ARQOS;
    output wire m_axi_gmem1_3_ARVALID;
    input wire m_axi_gmem1_3_ARREADY;
    input wire [63 : 0] m_axi_gmem1_3_RDATA;
    input wire [1 : 0] m_axi_gmem1_3_RRESP;
    input wire m_axi_gmem1_3_RLAST;
    input wire m_axi_gmem1_3_RVALID;
    output wire m_axi_gmem1_3_RREADY;
    output wire [63 : 0] m_axi_gmem1_4_AWADDR;
    output wire [7 : 0] m_axi_gmem1_4_AWLEN;
    output wire [2 : 0] m_axi_gmem1_4_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_4_AWBURST;
    output wire [1 : 0] m_axi_gmem1_4_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_4_AWREGION;
    output wire [3 : 0] m_axi_gmem1_4_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_4_AWPROT;
    output wire [3 : 0] m_axi_gmem1_4_AWQOS;
    output wire m_axi_gmem1_4_AWVALID;
    input wire m_axi_gmem1_4_AWREADY;
    output wire [63 : 0] m_axi_gmem1_4_WDATA;
    output wire [7 : 0] m_axi_gmem1_4_WSTRB;
    output wire m_axi_gmem1_4_WLAST;
    output wire m_axi_gmem1_4_WVALID;
    input wire m_axi_gmem1_4_WREADY;
    input wire [1 : 0] m_axi_gmem1_4_BRESP;
    input wire m_axi_gmem1_4_BVALID;
    output wire m_axi_gmem1_4_BREADY;
    output wire [63 : 0] m_axi_gmem1_4_ARADDR;
    output wire [7 : 0] m_axi_gmem1_4_ARLEN;
    output wire [2 : 0] m_axi_gmem1_4_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_4_ARBURST;
    output wire [1 : 0] m_axi_gmem1_4_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_4_ARREGION;
    output wire [3 : 0] m_axi_gmem1_4_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_4_ARPROT;
    output wire [3 : 0] m_axi_gmem1_4_ARQOS;
    output wire m_axi_gmem1_4_ARVALID;
    input wire m_axi_gmem1_4_ARREADY;
    input wire [63 : 0] m_axi_gmem1_4_RDATA;
    input wire [1 : 0] m_axi_gmem1_4_RRESP;
    input wire m_axi_gmem1_4_RLAST;
    input wire m_axi_gmem1_4_RVALID;
    output wire m_axi_gmem1_4_RREADY;
    output wire [63 : 0] m_axi_gmem1_5_AWADDR;
    output wire [7 : 0] m_axi_gmem1_5_AWLEN;
    output wire [2 : 0] m_axi_gmem1_5_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_5_AWBURST;
    output wire [1 : 0] m_axi_gmem1_5_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_5_AWREGION;
    output wire [3 : 0] m_axi_gmem1_5_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_5_AWPROT;
    output wire [3 : 0] m_axi_gmem1_5_AWQOS;
    output wire m_axi_gmem1_5_AWVALID;
    input wire m_axi_gmem1_5_AWREADY;
    output wire [63 : 0] m_axi_gmem1_5_WDATA;
    output wire [7 : 0] m_axi_gmem1_5_WSTRB;
    output wire m_axi_gmem1_5_WLAST;
    output wire m_axi_gmem1_5_WVALID;
    input wire m_axi_gmem1_5_WREADY;
    input wire [1 : 0] m_axi_gmem1_5_BRESP;
    input wire m_axi_gmem1_5_BVALID;
    output wire m_axi_gmem1_5_BREADY;
    output wire [63 : 0] m_axi_gmem1_5_ARADDR;
    output wire [7 : 0] m_axi_gmem1_5_ARLEN;
    output wire [2 : 0] m_axi_gmem1_5_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_5_ARBURST;
    output wire [1 : 0] m_axi_gmem1_5_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_5_ARREGION;
    output wire [3 : 0] m_axi_gmem1_5_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_5_ARPROT;
    output wire [3 : 0] m_axi_gmem1_5_ARQOS;
    output wire m_axi_gmem1_5_ARVALID;
    input wire m_axi_gmem1_5_ARREADY;
    input wire [63 : 0] m_axi_gmem1_5_RDATA;
    input wire [1 : 0] m_axi_gmem1_5_RRESP;
    input wire m_axi_gmem1_5_RLAST;
    input wire m_axi_gmem1_5_RVALID;
    output wire m_axi_gmem1_5_RREADY;
    output wire [63 : 0] m_axi_gmem1_6_AWADDR;
    output wire [7 : 0] m_axi_gmem1_6_AWLEN;
    output wire [2 : 0] m_axi_gmem1_6_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_6_AWBURST;
    output wire [1 : 0] m_axi_gmem1_6_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_6_AWREGION;
    output wire [3 : 0] m_axi_gmem1_6_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_6_AWPROT;
    output wire [3 : 0] m_axi_gmem1_6_AWQOS;
    output wire m_axi_gmem1_6_AWVALID;
    input wire m_axi_gmem1_6_AWREADY;
    output wire [63 : 0] m_axi_gmem1_6_WDATA;
    output wire [7 : 0] m_axi_gmem1_6_WSTRB;
    output wire m_axi_gmem1_6_WLAST;
    output wire m_axi_gmem1_6_WVALID;
    input wire m_axi_gmem1_6_WREADY;
    input wire [1 : 0] m_axi_gmem1_6_BRESP;
    input wire m_axi_gmem1_6_BVALID;
    output wire m_axi_gmem1_6_BREADY;
    output wire [63 : 0] m_axi_gmem1_6_ARADDR;
    output wire [7 : 0] m_axi_gmem1_6_ARLEN;
    output wire [2 : 0] m_axi_gmem1_6_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_6_ARBURST;
    output wire [1 : 0] m_axi_gmem1_6_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_6_ARREGION;
    output wire [3 : 0] m_axi_gmem1_6_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_6_ARPROT;
    output wire [3 : 0] m_axi_gmem1_6_ARQOS;
    output wire m_axi_gmem1_6_ARVALID;
    input wire m_axi_gmem1_6_ARREADY;
    input wire [63 : 0] m_axi_gmem1_6_RDATA;
    input wire [1 : 0] m_axi_gmem1_6_RRESP;
    input wire m_axi_gmem1_6_RLAST;
    input wire m_axi_gmem1_6_RVALID;
    output wire m_axi_gmem1_6_RREADY;
    output wire [63 : 0] m_axi_gmem1_7_AWADDR;
    output wire [7 : 0] m_axi_gmem1_7_AWLEN;
    output wire [2 : 0] m_axi_gmem1_7_AWSIZE;
    output wire [1 : 0] m_axi_gmem1_7_AWBURST;
    output wire [1 : 0] m_axi_gmem1_7_AWLOCK;
    output wire [3 : 0] m_axi_gmem1_7_AWREGION;
    output wire [3 : 0] m_axi_gmem1_7_AWCACHE;
    output wire [2 : 0] m_axi_gmem1_7_AWPROT;
    output wire [3 : 0] m_axi_gmem1_7_AWQOS;
    output wire m_axi_gmem1_7_AWVALID;
    input wire m_axi_gmem1_7_AWREADY;
    output wire [63 : 0] m_axi_gmem1_7_WDATA;
    output wire [7 : 0] m_axi_gmem1_7_WSTRB;
    output wire m_axi_gmem1_7_WLAST;
    output wire m_axi_gmem1_7_WVALID;
    input wire m_axi_gmem1_7_WREADY;
    input wire [1 : 0] m_axi_gmem1_7_BRESP;
    input wire m_axi_gmem1_7_BVALID;
    output wire m_axi_gmem1_7_BREADY;
    output wire [63 : 0] m_axi_gmem1_7_ARADDR;
    output wire [7 : 0] m_axi_gmem1_7_ARLEN;
    output wire [2 : 0] m_axi_gmem1_7_ARSIZE;
    output wire [1 : 0] m_axi_gmem1_7_ARBURST;
    output wire [1 : 0] m_axi_gmem1_7_ARLOCK;
    output wire [3 : 0] m_axi_gmem1_7_ARREGION;
    output wire [3 : 0] m_axi_gmem1_7_ARCACHE;
    output wire [2 : 0] m_axi_gmem1_7_ARPROT;
    output wire [3 : 0] m_axi_gmem1_7_ARQOS;
    output wire m_axi_gmem1_7_ARVALID;
    input wire m_axi_gmem1_7_ARREADY;
    input wire [63 : 0] m_axi_gmem1_7_RDATA;
    input wire [1 : 0] m_axi_gmem1_7_RRESP;
    input wire m_axi_gmem1_7_RLAST;
    input wire m_axi_gmem1_7_RVALID;
    output wire m_axi_gmem1_7_RREADY;
    output wire [63 : 0] m_axi_gmem2_0_AWADDR;
    output wire [7 : 0] m_axi_gmem2_0_AWLEN;
    output wire [2 : 0] m_axi_gmem2_0_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_0_AWBURST;
    output wire [1 : 0] m_axi_gmem2_0_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_0_AWREGION;
    output wire [3 : 0] m_axi_gmem2_0_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_0_AWPROT;
    output wire [3 : 0] m_axi_gmem2_0_AWQOS;
    output wire m_axi_gmem2_0_AWVALID;
    input wire m_axi_gmem2_0_AWREADY;
    output wire [63 : 0] m_axi_gmem2_0_WDATA;
    output wire [7 : 0] m_axi_gmem2_0_WSTRB;
    output wire m_axi_gmem2_0_WLAST;
    output wire m_axi_gmem2_0_WVALID;
    input wire m_axi_gmem2_0_WREADY;
    input wire [1 : 0] m_axi_gmem2_0_BRESP;
    input wire m_axi_gmem2_0_BVALID;
    output wire m_axi_gmem2_0_BREADY;
    output wire [63 : 0] m_axi_gmem2_0_ARADDR;
    output wire [7 : 0] m_axi_gmem2_0_ARLEN;
    output wire [2 : 0] m_axi_gmem2_0_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_0_ARBURST;
    output wire [1 : 0] m_axi_gmem2_0_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_0_ARREGION;
    output wire [3 : 0] m_axi_gmem2_0_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_0_ARPROT;
    output wire [3 : 0] m_axi_gmem2_0_ARQOS;
    output wire m_axi_gmem2_0_ARVALID;
    input wire m_axi_gmem2_0_ARREADY;
    input wire [63 : 0] m_axi_gmem2_0_RDATA;
    input wire [1 : 0] m_axi_gmem2_0_RRESP;
    input wire m_axi_gmem2_0_RLAST;
    input wire m_axi_gmem2_0_RVALID;
    output wire m_axi_gmem2_0_RREADY;
    output wire [63 : 0] m_axi_gmem2_1_AWADDR;
    output wire [7 : 0] m_axi_gmem2_1_AWLEN;
    output wire [2 : 0] m_axi_gmem2_1_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_1_AWBURST;
    output wire [1 : 0] m_axi_gmem2_1_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_1_AWREGION;
    output wire [3 : 0] m_axi_gmem2_1_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_1_AWPROT;
    output wire [3 : 0] m_axi_gmem2_1_AWQOS;
    output wire m_axi_gmem2_1_AWVALID;
    input wire m_axi_gmem2_1_AWREADY;
    output wire [63 : 0] m_axi_gmem2_1_WDATA;
    output wire [7 : 0] m_axi_gmem2_1_WSTRB;
    output wire m_axi_gmem2_1_WLAST;
    output wire m_axi_gmem2_1_WVALID;
    input wire m_axi_gmem2_1_WREADY;
    input wire [1 : 0] m_axi_gmem2_1_BRESP;
    input wire m_axi_gmem2_1_BVALID;
    output wire m_axi_gmem2_1_BREADY;
    output wire [63 : 0] m_axi_gmem2_1_ARADDR;
    output wire [7 : 0] m_axi_gmem2_1_ARLEN;
    output wire [2 : 0] m_axi_gmem2_1_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_1_ARBURST;
    output wire [1 : 0] m_axi_gmem2_1_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_1_ARREGION;
    output wire [3 : 0] m_axi_gmem2_1_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_1_ARPROT;
    output wire [3 : 0] m_axi_gmem2_1_ARQOS;
    output wire m_axi_gmem2_1_ARVALID;
    input wire m_axi_gmem2_1_ARREADY;
    input wire [63 : 0] m_axi_gmem2_1_RDATA;
    input wire [1 : 0] m_axi_gmem2_1_RRESP;
    input wire m_axi_gmem2_1_RLAST;
    input wire m_axi_gmem2_1_RVALID;
    output wire m_axi_gmem2_1_RREADY;
    output wire [63 : 0] m_axi_gmem2_2_AWADDR;
    output wire [7 : 0] m_axi_gmem2_2_AWLEN;
    output wire [2 : 0] m_axi_gmem2_2_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_2_AWBURST;
    output wire [1 : 0] m_axi_gmem2_2_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_2_AWREGION;
    output wire [3 : 0] m_axi_gmem2_2_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_2_AWPROT;
    output wire [3 : 0] m_axi_gmem2_2_AWQOS;
    output wire m_axi_gmem2_2_AWVALID;
    input wire m_axi_gmem2_2_AWREADY;
    output wire [63 : 0] m_axi_gmem2_2_WDATA;
    output wire [7 : 0] m_axi_gmem2_2_WSTRB;
    output wire m_axi_gmem2_2_WLAST;
    output wire m_axi_gmem2_2_WVALID;
    input wire m_axi_gmem2_2_WREADY;
    input wire [1 : 0] m_axi_gmem2_2_BRESP;
    input wire m_axi_gmem2_2_BVALID;
    output wire m_axi_gmem2_2_BREADY;
    output wire [63 : 0] m_axi_gmem2_2_ARADDR;
    output wire [7 : 0] m_axi_gmem2_2_ARLEN;
    output wire [2 : 0] m_axi_gmem2_2_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_2_ARBURST;
    output wire [1 : 0] m_axi_gmem2_2_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_2_ARREGION;
    output wire [3 : 0] m_axi_gmem2_2_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_2_ARPROT;
    output wire [3 : 0] m_axi_gmem2_2_ARQOS;
    output wire m_axi_gmem2_2_ARVALID;
    input wire m_axi_gmem2_2_ARREADY;
    input wire [63 : 0] m_axi_gmem2_2_RDATA;
    input wire [1 : 0] m_axi_gmem2_2_RRESP;
    input wire m_axi_gmem2_2_RLAST;
    input wire m_axi_gmem2_2_RVALID;
    output wire m_axi_gmem2_2_RREADY;
    output wire [63 : 0] m_axi_gmem2_3_AWADDR;
    output wire [7 : 0] m_axi_gmem2_3_AWLEN;
    output wire [2 : 0] m_axi_gmem2_3_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_3_AWBURST;
    output wire [1 : 0] m_axi_gmem2_3_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_3_AWREGION;
    output wire [3 : 0] m_axi_gmem2_3_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_3_AWPROT;
    output wire [3 : 0] m_axi_gmem2_3_AWQOS;
    output wire m_axi_gmem2_3_AWVALID;
    input wire m_axi_gmem2_3_AWREADY;
    output wire [63 : 0] m_axi_gmem2_3_WDATA;
    output wire [7 : 0] m_axi_gmem2_3_WSTRB;
    output wire m_axi_gmem2_3_WLAST;
    output wire m_axi_gmem2_3_WVALID;
    input wire m_axi_gmem2_3_WREADY;
    input wire [1 : 0] m_axi_gmem2_3_BRESP;
    input wire m_axi_gmem2_3_BVALID;
    output wire m_axi_gmem2_3_BREADY;
    output wire [63 : 0] m_axi_gmem2_3_ARADDR;
    output wire [7 : 0] m_axi_gmem2_3_ARLEN;
    output wire [2 : 0] m_axi_gmem2_3_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_3_ARBURST;
    output wire [1 : 0] m_axi_gmem2_3_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_3_ARREGION;
    output wire [3 : 0] m_axi_gmem2_3_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_3_ARPROT;
    output wire [3 : 0] m_axi_gmem2_3_ARQOS;
    output wire m_axi_gmem2_3_ARVALID;
    input wire m_axi_gmem2_3_ARREADY;
    input wire [63 : 0] m_axi_gmem2_3_RDATA;
    input wire [1 : 0] m_axi_gmem2_3_RRESP;
    input wire m_axi_gmem2_3_RLAST;
    input wire m_axi_gmem2_3_RVALID;
    output wire m_axi_gmem2_3_RREADY;
    output wire [63 : 0] m_axi_gmem2_4_AWADDR;
    output wire [7 : 0] m_axi_gmem2_4_AWLEN;
    output wire [2 : 0] m_axi_gmem2_4_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_4_AWBURST;
    output wire [1 : 0] m_axi_gmem2_4_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_4_AWREGION;
    output wire [3 : 0] m_axi_gmem2_4_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_4_AWPROT;
    output wire [3 : 0] m_axi_gmem2_4_AWQOS;
    output wire m_axi_gmem2_4_AWVALID;
    input wire m_axi_gmem2_4_AWREADY;
    output wire [63 : 0] m_axi_gmem2_4_WDATA;
    output wire [7 : 0] m_axi_gmem2_4_WSTRB;
    output wire m_axi_gmem2_4_WLAST;
    output wire m_axi_gmem2_4_WVALID;
    input wire m_axi_gmem2_4_WREADY;
    input wire [1 : 0] m_axi_gmem2_4_BRESP;
    input wire m_axi_gmem2_4_BVALID;
    output wire m_axi_gmem2_4_BREADY;
    output wire [63 : 0] m_axi_gmem2_4_ARADDR;
    output wire [7 : 0] m_axi_gmem2_4_ARLEN;
    output wire [2 : 0] m_axi_gmem2_4_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_4_ARBURST;
    output wire [1 : 0] m_axi_gmem2_4_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_4_ARREGION;
    output wire [3 : 0] m_axi_gmem2_4_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_4_ARPROT;
    output wire [3 : 0] m_axi_gmem2_4_ARQOS;
    output wire m_axi_gmem2_4_ARVALID;
    input wire m_axi_gmem2_4_ARREADY;
    input wire [63 : 0] m_axi_gmem2_4_RDATA;
    input wire [1 : 0] m_axi_gmem2_4_RRESP;
    input wire m_axi_gmem2_4_RLAST;
    input wire m_axi_gmem2_4_RVALID;
    output wire m_axi_gmem2_4_RREADY;
    output wire [63 : 0] m_axi_gmem2_5_AWADDR;
    output wire [7 : 0] m_axi_gmem2_5_AWLEN;
    output wire [2 : 0] m_axi_gmem2_5_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_5_AWBURST;
    output wire [1 : 0] m_axi_gmem2_5_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_5_AWREGION;
    output wire [3 : 0] m_axi_gmem2_5_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_5_AWPROT;
    output wire [3 : 0] m_axi_gmem2_5_AWQOS;
    output wire m_axi_gmem2_5_AWVALID;
    input wire m_axi_gmem2_5_AWREADY;
    output wire [63 : 0] m_axi_gmem2_5_WDATA;
    output wire [7 : 0] m_axi_gmem2_5_WSTRB;
    output wire m_axi_gmem2_5_WLAST;
    output wire m_axi_gmem2_5_WVALID;
    input wire m_axi_gmem2_5_WREADY;
    input wire [1 : 0] m_axi_gmem2_5_BRESP;
    input wire m_axi_gmem2_5_BVALID;
    output wire m_axi_gmem2_5_BREADY;
    output wire [63 : 0] m_axi_gmem2_5_ARADDR;
    output wire [7 : 0] m_axi_gmem2_5_ARLEN;
    output wire [2 : 0] m_axi_gmem2_5_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_5_ARBURST;
    output wire [1 : 0] m_axi_gmem2_5_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_5_ARREGION;
    output wire [3 : 0] m_axi_gmem2_5_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_5_ARPROT;
    output wire [3 : 0] m_axi_gmem2_5_ARQOS;
    output wire m_axi_gmem2_5_ARVALID;
    input wire m_axi_gmem2_5_ARREADY;
    input wire [63 : 0] m_axi_gmem2_5_RDATA;
    input wire [1 : 0] m_axi_gmem2_5_RRESP;
    input wire m_axi_gmem2_5_RLAST;
    input wire m_axi_gmem2_5_RVALID;
    output wire m_axi_gmem2_5_RREADY;
    output wire [63 : 0] m_axi_gmem2_6_AWADDR;
    output wire [7 : 0] m_axi_gmem2_6_AWLEN;
    output wire [2 : 0] m_axi_gmem2_6_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_6_AWBURST;
    output wire [1 : 0] m_axi_gmem2_6_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_6_AWREGION;
    output wire [3 : 0] m_axi_gmem2_6_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_6_AWPROT;
    output wire [3 : 0] m_axi_gmem2_6_AWQOS;
    output wire m_axi_gmem2_6_AWVALID;
    input wire m_axi_gmem2_6_AWREADY;
    output wire [63 : 0] m_axi_gmem2_6_WDATA;
    output wire [7 : 0] m_axi_gmem2_6_WSTRB;
    output wire m_axi_gmem2_6_WLAST;
    output wire m_axi_gmem2_6_WVALID;
    input wire m_axi_gmem2_6_WREADY;
    input wire [1 : 0] m_axi_gmem2_6_BRESP;
    input wire m_axi_gmem2_6_BVALID;
    output wire m_axi_gmem2_6_BREADY;
    output wire [63 : 0] m_axi_gmem2_6_ARADDR;
    output wire [7 : 0] m_axi_gmem2_6_ARLEN;
    output wire [2 : 0] m_axi_gmem2_6_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_6_ARBURST;
    output wire [1 : 0] m_axi_gmem2_6_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_6_ARREGION;
    output wire [3 : 0] m_axi_gmem2_6_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_6_ARPROT;
    output wire [3 : 0] m_axi_gmem2_6_ARQOS;
    output wire m_axi_gmem2_6_ARVALID;
    input wire m_axi_gmem2_6_ARREADY;
    input wire [63 : 0] m_axi_gmem2_6_RDATA;
    input wire [1 : 0] m_axi_gmem2_6_RRESP;
    input wire m_axi_gmem2_6_RLAST;
    input wire m_axi_gmem2_6_RVALID;
    output wire m_axi_gmem2_6_RREADY;
    output wire [63 : 0] m_axi_gmem2_7_AWADDR;
    output wire [7 : 0] m_axi_gmem2_7_AWLEN;
    output wire [2 : 0] m_axi_gmem2_7_AWSIZE;
    output wire [1 : 0] m_axi_gmem2_7_AWBURST;
    output wire [1 : 0] m_axi_gmem2_7_AWLOCK;
    output wire [3 : 0] m_axi_gmem2_7_AWREGION;
    output wire [3 : 0] m_axi_gmem2_7_AWCACHE;
    output wire [2 : 0] m_axi_gmem2_7_AWPROT;
    output wire [3 : 0] m_axi_gmem2_7_AWQOS;
    output wire m_axi_gmem2_7_AWVALID;
    input wire m_axi_gmem2_7_AWREADY;
    output wire [63 : 0] m_axi_gmem2_7_WDATA;
    output wire [7 : 0] m_axi_gmem2_7_WSTRB;
    output wire m_axi_gmem2_7_WLAST;
    output wire m_axi_gmem2_7_WVALID;
    input wire m_axi_gmem2_7_WREADY;
    input wire [1 : 0] m_axi_gmem2_7_BRESP;
    input wire m_axi_gmem2_7_BVALID;
    output wire m_axi_gmem2_7_BREADY;
    output wire [63 : 0] m_axi_gmem2_7_ARADDR;
    output wire [7 : 0] m_axi_gmem2_7_ARLEN;
    output wire [2 : 0] m_axi_gmem2_7_ARSIZE;
    output wire [1 : 0] m_axi_gmem2_7_ARBURST;
    output wire [1 : 0] m_axi_gmem2_7_ARLOCK;
    output wire [3 : 0] m_axi_gmem2_7_ARREGION;
    output wire [3 : 0] m_axi_gmem2_7_ARCACHE;
    output wire [2 : 0] m_axi_gmem2_7_ARPROT;
    output wire [3 : 0] m_axi_gmem2_7_ARQOS;
    output wire m_axi_gmem2_7_ARVALID;
    input wire m_axi_gmem2_7_ARREADY;
    input wire [63 : 0] m_axi_gmem2_7_RDATA;
    input wire [1 : 0] m_axi_gmem2_7_RRESP;
    input wire m_axi_gmem2_7_RLAST;
    input wire m_axi_gmem2_7_RVALID;
    output wire m_axi_gmem2_7_RREADY;

    gqeJoin_1 gqeJoin_1_0     (
        .stall_start_ext        ( stall_start_ext        ) , // output wire stall_start_ext
        .stall_done_ext         ( stall_done_ext         ) , // output wire stall_done_ext
        .stall_start_str        ( stall_start_str        ) , // output wire stall_start_str
        .stall_done_str         ( stall_done_str         ) , // output wire stall_done_str
        .stall_start_int        ( stall_start_int        ) , // output wire stall_start_int
        .stall_done_int         ( stall_done_int         ) , // output wire stall_done_int
        .s_axi_control_AWADDR   ( s_axi_control_AWADDR   ) , // input wire [7 : 0] s_axi_control_AWADDR
        .s_axi_control_AWVALID  ( s_axi_control_AWVALID  ) , // input wire s_axi_control_AWVALID
        .s_axi_control_AWREADY  ( s_axi_control_AWREADY  ) , // output wire s_axi_control_AWREADY
        .s_axi_control_WDATA    ( s_axi_control_WDATA    ) , // input wire [31 : 0] s_axi_control_WDATA
        .s_axi_control_WSTRB    ( s_axi_control_WSTRB    ) , // input wire [3 : 0] s_axi_control_WSTRB
        .s_axi_control_WVALID   ( s_axi_control_WVALID   ) , // input wire s_axi_control_WVALID
        .s_axi_control_WREADY   ( s_axi_control_WREADY   ) , // output wire s_axi_control_WREADY
        .s_axi_control_BRESP    ( s_axi_control_BRESP    ) , // output wire [1 : 0] s_axi_control_BRESP
        .s_axi_control_BVALID   ( s_axi_control_BVALID   ) , // output wire s_axi_control_BVALID
        .s_axi_control_BREADY   ( s_axi_control_BREADY   ) , // input wire s_axi_control_BREADY
        .s_axi_control_ARADDR   ( s_axi_control_ARADDR   ) , // input wire [7 : 0] s_axi_control_ARADDR
        .s_axi_control_ARVALID  ( s_axi_control_ARVALID  ) , // input wire s_axi_control_ARVALID
        .s_axi_control_ARREADY  ( s_axi_control_ARREADY  ) , // output wire s_axi_control_ARREADY
        .s_axi_control_RDATA    ( s_axi_control_RDATA    ) , // output wire [31 : 0] s_axi_control_RDATA
        .s_axi_control_RRESP    ( s_axi_control_RRESP    ) , // output wire [1 : 0] s_axi_control_RRESP
        .s_axi_control_RVALID   ( s_axi_control_RVALID   ) , // output wire s_axi_control_RVALID
        .s_axi_control_RREADY   ( s_axi_control_RREADY   ) , // input wire s_axi_control_RREADY
        .ap_clk                 ( ap_clk                 ) , // input wire ap_clk
        .ap_rst_n               ( ap_rst_n               ) , // input wire ap_rst_n
        .event_done             ( event_done             ) , // output wire event_done
        .interrupt              ( interrupt              ) , // output wire interrupt
        .event_start            ( event_start            ) , // output wire event_start
        .m_axi_gmem0_0_AWADDR   ( m_axi_gmem0_0_AWADDR   ) , // output wire [63 : 0] m_axi_gmem0_0_AWADDR
        .m_axi_gmem0_0_AWLEN    ( m_axi_gmem0_0_AWLEN    ) , // output wire [7 : 0] m_axi_gmem0_0_AWLEN
        .m_axi_gmem0_0_AWSIZE   ( m_axi_gmem0_0_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem0_0_AWSIZE
        .m_axi_gmem0_0_AWBURST  ( m_axi_gmem0_0_AWBURST  ) , // output wire [1 : 0] m_axi_gmem0_0_AWBURST
        .m_axi_gmem0_0_AWLOCK   ( m_axi_gmem0_0_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem0_0_AWLOCK
        .m_axi_gmem0_0_AWREGION ( m_axi_gmem0_0_AWREGION ) , // output wire [3 : 0] m_axi_gmem0_0_AWREGION
        .m_axi_gmem0_0_AWCACHE  ( m_axi_gmem0_0_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem0_0_AWCACHE
        .m_axi_gmem0_0_AWPROT   ( m_axi_gmem0_0_AWPROT   ) , // output wire [2 : 0] m_axi_gmem0_0_AWPROT
        .m_axi_gmem0_0_AWQOS    ( m_axi_gmem0_0_AWQOS    ) , // output wire [3 : 0] m_axi_gmem0_0_AWQOS
        .m_axi_gmem0_0_AWVALID  ( m_axi_gmem0_0_AWVALID  ) , // output wire m_axi_gmem0_0_AWVALID
        .m_axi_gmem0_0_AWREADY  ( m_axi_gmem0_0_AWREADY  ) , // input wire m_axi_gmem0_0_AWREADY
        .m_axi_gmem0_0_WDATA    ( m_axi_gmem0_0_WDATA    ) , // output wire [511 : 0] m_axi_gmem0_0_WDATA
        .m_axi_gmem0_0_WSTRB    ( m_axi_gmem0_0_WSTRB    ) , // output wire [63 : 0] m_axi_gmem0_0_WSTRB
        .m_axi_gmem0_0_WLAST    ( m_axi_gmem0_0_WLAST    ) , // output wire m_axi_gmem0_0_WLAST
        .m_axi_gmem0_0_WVALID   ( m_axi_gmem0_0_WVALID   ) , // output wire m_axi_gmem0_0_WVALID
        .m_axi_gmem0_0_WREADY   ( m_axi_gmem0_0_WREADY   ) , // input wire m_axi_gmem0_0_WREADY
        .m_axi_gmem0_0_BRESP    ( m_axi_gmem0_0_BRESP    ) , // input wire [1 : 0] m_axi_gmem0_0_BRESP
        .m_axi_gmem0_0_BVALID   ( m_axi_gmem0_0_BVALID   ) , // input wire m_axi_gmem0_0_BVALID
        .m_axi_gmem0_0_BREADY   ( m_axi_gmem0_0_BREADY   ) , // output wire m_axi_gmem0_0_BREADY
        .m_axi_gmem0_0_ARADDR   ( m_axi_gmem0_0_ARADDR   ) , // output wire [63 : 0] m_axi_gmem0_0_ARADDR
        .m_axi_gmem0_0_ARLEN    ( m_axi_gmem0_0_ARLEN    ) , // output wire [7 : 0] m_axi_gmem0_0_ARLEN
        .m_axi_gmem0_0_ARSIZE   ( m_axi_gmem0_0_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem0_0_ARSIZE
        .m_axi_gmem0_0_ARBURST  ( m_axi_gmem0_0_ARBURST  ) , // output wire [1 : 0] m_axi_gmem0_0_ARBURST
        .m_axi_gmem0_0_ARLOCK   ( m_axi_gmem0_0_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem0_0_ARLOCK
        .m_axi_gmem0_0_ARREGION ( m_axi_gmem0_0_ARREGION ) , // output wire [3 : 0] m_axi_gmem0_0_ARREGION
        .m_axi_gmem0_0_ARCACHE  ( m_axi_gmem0_0_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem0_0_ARCACHE
        .m_axi_gmem0_0_ARPROT   ( m_axi_gmem0_0_ARPROT   ) , // output wire [2 : 0] m_axi_gmem0_0_ARPROT
        .m_axi_gmem0_0_ARQOS    ( m_axi_gmem0_0_ARQOS    ) , // output wire [3 : 0] m_axi_gmem0_0_ARQOS
        .m_axi_gmem0_0_ARVALID  ( m_axi_gmem0_0_ARVALID  ) , // output wire m_axi_gmem0_0_ARVALID
        .m_axi_gmem0_0_ARREADY  ( m_axi_gmem0_0_ARREADY  ) , // input wire m_axi_gmem0_0_ARREADY
        .m_axi_gmem0_0_RDATA    ( m_axi_gmem0_0_RDATA    ) , // input wire [511 : 0] m_axi_gmem0_0_RDATA
        .m_axi_gmem0_0_RRESP    ( m_axi_gmem0_0_RRESP    ) , // input wire [1 : 0] m_axi_gmem0_0_RRESP
        .m_axi_gmem0_0_RLAST    ( m_axi_gmem0_0_RLAST    ) , // input wire m_axi_gmem0_0_RLAST
        .m_axi_gmem0_0_RVALID   ( m_axi_gmem0_0_RVALID   ) , // input wire m_axi_gmem0_0_RVALID
        .m_axi_gmem0_0_RREADY   ( m_axi_gmem0_0_RREADY   ) , // output wire m_axi_gmem0_0_RREADY
        .m_axi_gmem0_1_AWADDR   ( m_axi_gmem0_1_AWADDR   ) , // output wire [63 : 0] m_axi_gmem0_1_AWADDR
        .m_axi_gmem0_1_AWLEN    ( m_axi_gmem0_1_AWLEN    ) , // output wire [7 : 0] m_axi_gmem0_1_AWLEN
        .m_axi_gmem0_1_AWSIZE   ( m_axi_gmem0_1_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem0_1_AWSIZE
        .m_axi_gmem0_1_AWBURST  ( m_axi_gmem0_1_AWBURST  ) , // output wire [1 : 0] m_axi_gmem0_1_AWBURST
        .m_axi_gmem0_1_AWLOCK   ( m_axi_gmem0_1_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem0_1_AWLOCK
        .m_axi_gmem0_1_AWREGION ( m_axi_gmem0_1_AWREGION ) , // output wire [3 : 0] m_axi_gmem0_1_AWREGION
        .m_axi_gmem0_1_AWCACHE  ( m_axi_gmem0_1_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem0_1_AWCACHE
        .m_axi_gmem0_1_AWPROT   ( m_axi_gmem0_1_AWPROT   ) , // output wire [2 : 0] m_axi_gmem0_1_AWPROT
        .m_axi_gmem0_1_AWQOS    ( m_axi_gmem0_1_AWQOS    ) , // output wire [3 : 0] m_axi_gmem0_1_AWQOS
        .m_axi_gmem0_1_AWVALID  ( m_axi_gmem0_1_AWVALID  ) , // output wire m_axi_gmem0_1_AWVALID
        .m_axi_gmem0_1_AWREADY  ( m_axi_gmem0_1_AWREADY  ) , // input wire m_axi_gmem0_1_AWREADY
        .m_axi_gmem0_1_WDATA    ( m_axi_gmem0_1_WDATA    ) , // output wire [511 : 0] m_axi_gmem0_1_WDATA
        .m_axi_gmem0_1_WSTRB    ( m_axi_gmem0_1_WSTRB    ) , // output wire [63 : 0] m_axi_gmem0_1_WSTRB
        .m_axi_gmem0_1_WLAST    ( m_axi_gmem0_1_WLAST    ) , // output wire m_axi_gmem0_1_WLAST
        .m_axi_gmem0_1_WVALID   ( m_axi_gmem0_1_WVALID   ) , // output wire m_axi_gmem0_1_WVALID
        .m_axi_gmem0_1_WREADY   ( m_axi_gmem0_1_WREADY   ) , // input wire m_axi_gmem0_1_WREADY
        .m_axi_gmem0_1_BRESP    ( m_axi_gmem0_1_BRESP    ) , // input wire [1 : 0] m_axi_gmem0_1_BRESP
        .m_axi_gmem0_1_BVALID   ( m_axi_gmem0_1_BVALID   ) , // input wire m_axi_gmem0_1_BVALID
        .m_axi_gmem0_1_BREADY   ( m_axi_gmem0_1_BREADY   ) , // output wire m_axi_gmem0_1_BREADY
        .m_axi_gmem0_1_ARADDR   ( m_axi_gmem0_1_ARADDR   ) , // output wire [63 : 0] m_axi_gmem0_1_ARADDR
        .m_axi_gmem0_1_ARLEN    ( m_axi_gmem0_1_ARLEN    ) , // output wire [7 : 0] m_axi_gmem0_1_ARLEN
        .m_axi_gmem0_1_ARSIZE   ( m_axi_gmem0_1_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem0_1_ARSIZE
        .m_axi_gmem0_1_ARBURST  ( m_axi_gmem0_1_ARBURST  ) , // output wire [1 : 0] m_axi_gmem0_1_ARBURST
        .m_axi_gmem0_1_ARLOCK   ( m_axi_gmem0_1_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem0_1_ARLOCK
        .m_axi_gmem0_1_ARREGION ( m_axi_gmem0_1_ARREGION ) , // output wire [3 : 0] m_axi_gmem0_1_ARREGION
        .m_axi_gmem0_1_ARCACHE  ( m_axi_gmem0_1_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem0_1_ARCACHE
        .m_axi_gmem0_1_ARPROT   ( m_axi_gmem0_1_ARPROT   ) , // output wire [2 : 0] m_axi_gmem0_1_ARPROT
        .m_axi_gmem0_1_ARQOS    ( m_axi_gmem0_1_ARQOS    ) , // output wire [3 : 0] m_axi_gmem0_1_ARQOS
        .m_axi_gmem0_1_ARVALID  ( m_axi_gmem0_1_ARVALID  ) , // output wire m_axi_gmem0_1_ARVALID
        .m_axi_gmem0_1_ARREADY  ( m_axi_gmem0_1_ARREADY  ) , // input wire m_axi_gmem0_1_ARREADY
        .m_axi_gmem0_1_RDATA    ( m_axi_gmem0_1_RDATA    ) , // input wire [511 : 0] m_axi_gmem0_1_RDATA
        .m_axi_gmem0_1_RRESP    ( m_axi_gmem0_1_RRESP    ) , // input wire [1 : 0] m_axi_gmem0_1_RRESP
        .m_axi_gmem0_1_RLAST    ( m_axi_gmem0_1_RLAST    ) , // input wire m_axi_gmem0_1_RLAST
        .m_axi_gmem0_1_RVALID   ( m_axi_gmem0_1_RVALID   ) , // input wire m_axi_gmem0_1_RVALID
        .m_axi_gmem0_1_RREADY   ( m_axi_gmem0_1_RREADY   ) , // output wire m_axi_gmem0_1_RREADY
        .m_axi_gmem0_2_AWADDR   ( m_axi_gmem0_2_AWADDR   ) , // output wire [63 : 0] m_axi_gmem0_2_AWADDR
        .m_axi_gmem0_2_AWLEN    ( m_axi_gmem0_2_AWLEN    ) , // output wire [7 : 0] m_axi_gmem0_2_AWLEN
        .m_axi_gmem0_2_AWSIZE   ( m_axi_gmem0_2_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem0_2_AWSIZE
        .m_axi_gmem0_2_AWBURST  ( m_axi_gmem0_2_AWBURST  ) , // output wire [1 : 0] m_axi_gmem0_2_AWBURST
        .m_axi_gmem0_2_AWLOCK   ( m_axi_gmem0_2_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem0_2_AWLOCK
        .m_axi_gmem0_2_AWREGION ( m_axi_gmem0_2_AWREGION ) , // output wire [3 : 0] m_axi_gmem0_2_AWREGION
        .m_axi_gmem0_2_AWCACHE  ( m_axi_gmem0_2_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem0_2_AWCACHE
        .m_axi_gmem0_2_AWPROT   ( m_axi_gmem0_2_AWPROT   ) , // output wire [2 : 0] m_axi_gmem0_2_AWPROT
        .m_axi_gmem0_2_AWQOS    ( m_axi_gmem0_2_AWQOS    ) , // output wire [3 : 0] m_axi_gmem0_2_AWQOS
        .m_axi_gmem0_2_AWVALID  ( m_axi_gmem0_2_AWVALID  ) , // output wire m_axi_gmem0_2_AWVALID
        .m_axi_gmem0_2_AWREADY  ( m_axi_gmem0_2_AWREADY  ) , // input wire m_axi_gmem0_2_AWREADY
        .m_axi_gmem0_2_WDATA    ( m_axi_gmem0_2_WDATA    ) , // output wire [511 : 0] m_axi_gmem0_2_WDATA
        .m_axi_gmem0_2_WSTRB    ( m_axi_gmem0_2_WSTRB    ) , // output wire [63 : 0] m_axi_gmem0_2_WSTRB
        .m_axi_gmem0_2_WLAST    ( m_axi_gmem0_2_WLAST    ) , // output wire m_axi_gmem0_2_WLAST
        .m_axi_gmem0_2_WVALID   ( m_axi_gmem0_2_WVALID   ) , // output wire m_axi_gmem0_2_WVALID
        .m_axi_gmem0_2_WREADY   ( m_axi_gmem0_2_WREADY   ) , // input wire m_axi_gmem0_2_WREADY
        .m_axi_gmem0_2_BRESP    ( m_axi_gmem0_2_BRESP    ) , // input wire [1 : 0] m_axi_gmem0_2_BRESP
        .m_axi_gmem0_2_BVALID   ( m_axi_gmem0_2_BVALID   ) , // input wire m_axi_gmem0_2_BVALID
        .m_axi_gmem0_2_BREADY   ( m_axi_gmem0_2_BREADY   ) , // output wire m_axi_gmem0_2_BREADY
        .m_axi_gmem0_2_ARADDR   ( m_axi_gmem0_2_ARADDR   ) , // output wire [63 : 0] m_axi_gmem0_2_ARADDR
        .m_axi_gmem0_2_ARLEN    ( m_axi_gmem0_2_ARLEN    ) , // output wire [7 : 0] m_axi_gmem0_2_ARLEN
        .m_axi_gmem0_2_ARSIZE   ( m_axi_gmem0_2_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem0_2_ARSIZE
        .m_axi_gmem0_2_ARBURST  ( m_axi_gmem0_2_ARBURST  ) , // output wire [1 : 0] m_axi_gmem0_2_ARBURST
        .m_axi_gmem0_2_ARLOCK   ( m_axi_gmem0_2_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem0_2_ARLOCK
        .m_axi_gmem0_2_ARREGION ( m_axi_gmem0_2_ARREGION ) , // output wire [3 : 0] m_axi_gmem0_2_ARREGION
        .m_axi_gmem0_2_ARCACHE  ( m_axi_gmem0_2_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem0_2_ARCACHE
        .m_axi_gmem0_2_ARPROT   ( m_axi_gmem0_2_ARPROT   ) , // output wire [2 : 0] m_axi_gmem0_2_ARPROT
        .m_axi_gmem0_2_ARQOS    ( m_axi_gmem0_2_ARQOS    ) , // output wire [3 : 0] m_axi_gmem0_2_ARQOS
        .m_axi_gmem0_2_ARVALID  ( m_axi_gmem0_2_ARVALID  ) , // output wire m_axi_gmem0_2_ARVALID
        .m_axi_gmem0_2_ARREADY  ( m_axi_gmem0_2_ARREADY  ) , // input wire m_axi_gmem0_2_ARREADY
        .m_axi_gmem0_2_RDATA    ( m_axi_gmem0_2_RDATA    ) , // input wire [511 : 0] m_axi_gmem0_2_RDATA
        .m_axi_gmem0_2_RRESP    ( m_axi_gmem0_2_RRESP    ) , // input wire [1 : 0] m_axi_gmem0_2_RRESP
        .m_axi_gmem0_2_RLAST    ( m_axi_gmem0_2_RLAST    ) , // input wire m_axi_gmem0_2_RLAST
        .m_axi_gmem0_2_RVALID   ( m_axi_gmem0_2_RVALID   ) , // input wire m_axi_gmem0_2_RVALID
        .m_axi_gmem0_2_RREADY   ( m_axi_gmem0_2_RREADY   ) , // output wire m_axi_gmem0_2_RREADY
        .m_axi_gmem0_3_AWADDR   ( m_axi_gmem0_3_AWADDR   ) , // output wire [63 : 0] m_axi_gmem0_3_AWADDR
        .m_axi_gmem0_3_AWLEN    ( m_axi_gmem0_3_AWLEN    ) , // output wire [7 : 0] m_axi_gmem0_3_AWLEN
        .m_axi_gmem0_3_AWSIZE   ( m_axi_gmem0_3_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem0_3_AWSIZE
        .m_axi_gmem0_3_AWBURST  ( m_axi_gmem0_3_AWBURST  ) , // output wire [1 : 0] m_axi_gmem0_3_AWBURST
        .m_axi_gmem0_3_AWLOCK   ( m_axi_gmem0_3_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem0_3_AWLOCK
        .m_axi_gmem0_3_AWREGION ( m_axi_gmem0_3_AWREGION ) , // output wire [3 : 0] m_axi_gmem0_3_AWREGION
        .m_axi_gmem0_3_AWCACHE  ( m_axi_gmem0_3_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem0_3_AWCACHE
        .m_axi_gmem0_3_AWPROT   ( m_axi_gmem0_3_AWPROT   ) , // output wire [2 : 0] m_axi_gmem0_3_AWPROT
        .m_axi_gmem0_3_AWQOS    ( m_axi_gmem0_3_AWQOS    ) , // output wire [3 : 0] m_axi_gmem0_3_AWQOS
        .m_axi_gmem0_3_AWVALID  ( m_axi_gmem0_3_AWVALID  ) , // output wire m_axi_gmem0_3_AWVALID
        .m_axi_gmem0_3_AWREADY  ( m_axi_gmem0_3_AWREADY  ) , // input wire m_axi_gmem0_3_AWREADY
        .m_axi_gmem0_3_WDATA    ( m_axi_gmem0_3_WDATA    ) , // output wire [511 : 0] m_axi_gmem0_3_WDATA
        .m_axi_gmem0_3_WSTRB    ( m_axi_gmem0_3_WSTRB    ) , // output wire [63 : 0] m_axi_gmem0_3_WSTRB
        .m_axi_gmem0_3_WLAST    ( m_axi_gmem0_3_WLAST    ) , // output wire m_axi_gmem0_3_WLAST
        .m_axi_gmem0_3_WVALID   ( m_axi_gmem0_3_WVALID   ) , // output wire m_axi_gmem0_3_WVALID
        .m_axi_gmem0_3_WREADY   ( m_axi_gmem0_3_WREADY   ) , // input wire m_axi_gmem0_3_WREADY
        .m_axi_gmem0_3_BRESP    ( m_axi_gmem0_3_BRESP    ) , // input wire [1 : 0] m_axi_gmem0_3_BRESP
        .m_axi_gmem0_3_BVALID   ( m_axi_gmem0_3_BVALID   ) , // input wire m_axi_gmem0_3_BVALID
        .m_axi_gmem0_3_BREADY   ( m_axi_gmem0_3_BREADY   ) , // output wire m_axi_gmem0_3_BREADY
        .m_axi_gmem0_3_ARADDR   ( m_axi_gmem0_3_ARADDR   ) , // output wire [63 : 0] m_axi_gmem0_3_ARADDR
        .m_axi_gmem0_3_ARLEN    ( m_axi_gmem0_3_ARLEN    ) , // output wire [7 : 0] m_axi_gmem0_3_ARLEN
        .m_axi_gmem0_3_ARSIZE   ( m_axi_gmem0_3_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem0_3_ARSIZE
        .m_axi_gmem0_3_ARBURST  ( m_axi_gmem0_3_ARBURST  ) , // output wire [1 : 0] m_axi_gmem0_3_ARBURST
        .m_axi_gmem0_3_ARLOCK   ( m_axi_gmem0_3_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem0_3_ARLOCK
        .m_axi_gmem0_3_ARREGION ( m_axi_gmem0_3_ARREGION ) , // output wire [3 : 0] m_axi_gmem0_3_ARREGION
        .m_axi_gmem0_3_ARCACHE  ( m_axi_gmem0_3_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem0_3_ARCACHE
        .m_axi_gmem0_3_ARPROT   ( m_axi_gmem0_3_ARPROT   ) , // output wire [2 : 0] m_axi_gmem0_3_ARPROT
        .m_axi_gmem0_3_ARQOS    ( m_axi_gmem0_3_ARQOS    ) , // output wire [3 : 0] m_axi_gmem0_3_ARQOS
        .m_axi_gmem0_3_ARVALID  ( m_axi_gmem0_3_ARVALID  ) , // output wire m_axi_gmem0_3_ARVALID
        .m_axi_gmem0_3_ARREADY  ( m_axi_gmem0_3_ARREADY  ) , // input wire m_axi_gmem0_3_ARREADY
        .m_axi_gmem0_3_RDATA    ( m_axi_gmem0_3_RDATA    ) , // input wire [511 : 0] m_axi_gmem0_3_RDATA
        .m_axi_gmem0_3_RRESP    ( m_axi_gmem0_3_RRESP    ) , // input wire [1 : 0] m_axi_gmem0_3_RRESP
        .m_axi_gmem0_3_RLAST    ( m_axi_gmem0_3_RLAST    ) , // input wire m_axi_gmem0_3_RLAST
        .m_axi_gmem0_3_RVALID   ( m_axi_gmem0_3_RVALID   ) , // input wire m_axi_gmem0_3_RVALID
        .m_axi_gmem0_3_RREADY   ( m_axi_gmem0_3_RREADY   ) , // output wire m_axi_gmem0_3_RREADY
        .m_axi_gmem1_0_AWADDR   ( m_axi_gmem1_0_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_0_AWADDR
        .m_axi_gmem1_0_AWLEN    ( m_axi_gmem1_0_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_0_AWLEN
        .m_axi_gmem1_0_AWSIZE   ( m_axi_gmem1_0_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_0_AWSIZE
        .m_axi_gmem1_0_AWBURST  ( m_axi_gmem1_0_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_0_AWBURST
        .m_axi_gmem1_0_AWLOCK   ( m_axi_gmem1_0_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_0_AWLOCK
        .m_axi_gmem1_0_AWREGION ( m_axi_gmem1_0_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_0_AWREGION
        .m_axi_gmem1_0_AWCACHE  ( m_axi_gmem1_0_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_0_AWCACHE
        .m_axi_gmem1_0_AWPROT   ( m_axi_gmem1_0_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_0_AWPROT
        .m_axi_gmem1_0_AWQOS    ( m_axi_gmem1_0_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_0_AWQOS
        .m_axi_gmem1_0_AWVALID  ( m_axi_gmem1_0_AWVALID  ) , // output wire m_axi_gmem1_0_AWVALID
        .m_axi_gmem1_0_AWREADY  ( m_axi_gmem1_0_AWREADY  ) , // input wire m_axi_gmem1_0_AWREADY
        .m_axi_gmem1_0_WDATA    ( m_axi_gmem1_0_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_0_WDATA
        .m_axi_gmem1_0_WSTRB    ( m_axi_gmem1_0_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_0_WSTRB
        .m_axi_gmem1_0_WLAST    ( m_axi_gmem1_0_WLAST    ) , // output wire m_axi_gmem1_0_WLAST
        .m_axi_gmem1_0_WVALID   ( m_axi_gmem1_0_WVALID   ) , // output wire m_axi_gmem1_0_WVALID
        .m_axi_gmem1_0_WREADY   ( m_axi_gmem1_0_WREADY   ) , // input wire m_axi_gmem1_0_WREADY
        .m_axi_gmem1_0_BRESP    ( m_axi_gmem1_0_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_0_BRESP
        .m_axi_gmem1_0_BVALID   ( m_axi_gmem1_0_BVALID   ) , // input wire m_axi_gmem1_0_BVALID
        .m_axi_gmem1_0_BREADY   ( m_axi_gmem1_0_BREADY   ) , // output wire m_axi_gmem1_0_BREADY
        .m_axi_gmem1_0_ARADDR   ( m_axi_gmem1_0_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_0_ARADDR
        .m_axi_gmem1_0_ARLEN    ( m_axi_gmem1_0_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_0_ARLEN
        .m_axi_gmem1_0_ARSIZE   ( m_axi_gmem1_0_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_0_ARSIZE
        .m_axi_gmem1_0_ARBURST  ( m_axi_gmem1_0_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_0_ARBURST
        .m_axi_gmem1_0_ARLOCK   ( m_axi_gmem1_0_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_0_ARLOCK
        .m_axi_gmem1_0_ARREGION ( m_axi_gmem1_0_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_0_ARREGION
        .m_axi_gmem1_0_ARCACHE  ( m_axi_gmem1_0_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_0_ARCACHE
        .m_axi_gmem1_0_ARPROT   ( m_axi_gmem1_0_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_0_ARPROT
        .m_axi_gmem1_0_ARQOS    ( m_axi_gmem1_0_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_0_ARQOS
        .m_axi_gmem1_0_ARVALID  ( m_axi_gmem1_0_ARVALID  ) , // output wire m_axi_gmem1_0_ARVALID
        .m_axi_gmem1_0_ARREADY  ( m_axi_gmem1_0_ARREADY  ) , // input wire m_axi_gmem1_0_ARREADY
        .m_axi_gmem1_0_RDATA    ( m_axi_gmem1_0_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_0_RDATA
        .m_axi_gmem1_0_RRESP    ( m_axi_gmem1_0_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_0_RRESP
        .m_axi_gmem1_0_RLAST    ( m_axi_gmem1_0_RLAST    ) , // input wire m_axi_gmem1_0_RLAST
        .m_axi_gmem1_0_RVALID   ( m_axi_gmem1_0_RVALID   ) , // input wire m_axi_gmem1_0_RVALID
        .m_axi_gmem1_0_RREADY   ( m_axi_gmem1_0_RREADY   ) , // output wire m_axi_gmem1_0_RREADY
        .m_axi_gmem1_1_AWADDR   ( m_axi_gmem1_1_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_1_AWADDR
        .m_axi_gmem1_1_AWLEN    ( m_axi_gmem1_1_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_1_AWLEN
        .m_axi_gmem1_1_AWSIZE   ( m_axi_gmem1_1_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_1_AWSIZE
        .m_axi_gmem1_1_AWBURST  ( m_axi_gmem1_1_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_1_AWBURST
        .m_axi_gmem1_1_AWLOCK   ( m_axi_gmem1_1_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_1_AWLOCK
        .m_axi_gmem1_1_AWREGION ( m_axi_gmem1_1_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_1_AWREGION
        .m_axi_gmem1_1_AWCACHE  ( m_axi_gmem1_1_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_1_AWCACHE
        .m_axi_gmem1_1_AWPROT   ( m_axi_gmem1_1_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_1_AWPROT
        .m_axi_gmem1_1_AWQOS    ( m_axi_gmem1_1_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_1_AWQOS
        .m_axi_gmem1_1_AWVALID  ( m_axi_gmem1_1_AWVALID  ) , // output wire m_axi_gmem1_1_AWVALID
        .m_axi_gmem1_1_AWREADY  ( m_axi_gmem1_1_AWREADY  ) , // input wire m_axi_gmem1_1_AWREADY
        .m_axi_gmem1_1_WDATA    ( m_axi_gmem1_1_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_1_WDATA
        .m_axi_gmem1_1_WSTRB    ( m_axi_gmem1_1_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_1_WSTRB
        .m_axi_gmem1_1_WLAST    ( m_axi_gmem1_1_WLAST    ) , // output wire m_axi_gmem1_1_WLAST
        .m_axi_gmem1_1_WVALID   ( m_axi_gmem1_1_WVALID   ) , // output wire m_axi_gmem1_1_WVALID
        .m_axi_gmem1_1_WREADY   ( m_axi_gmem1_1_WREADY   ) , // input wire m_axi_gmem1_1_WREADY
        .m_axi_gmem1_1_BRESP    ( m_axi_gmem1_1_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_1_BRESP
        .m_axi_gmem1_1_BVALID   ( m_axi_gmem1_1_BVALID   ) , // input wire m_axi_gmem1_1_BVALID
        .m_axi_gmem1_1_BREADY   ( m_axi_gmem1_1_BREADY   ) , // output wire m_axi_gmem1_1_BREADY
        .m_axi_gmem1_1_ARADDR   ( m_axi_gmem1_1_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_1_ARADDR
        .m_axi_gmem1_1_ARLEN    ( m_axi_gmem1_1_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_1_ARLEN
        .m_axi_gmem1_1_ARSIZE   ( m_axi_gmem1_1_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_1_ARSIZE
        .m_axi_gmem1_1_ARBURST  ( m_axi_gmem1_1_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_1_ARBURST
        .m_axi_gmem1_1_ARLOCK   ( m_axi_gmem1_1_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_1_ARLOCK
        .m_axi_gmem1_1_ARREGION ( m_axi_gmem1_1_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_1_ARREGION
        .m_axi_gmem1_1_ARCACHE  ( m_axi_gmem1_1_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_1_ARCACHE
        .m_axi_gmem1_1_ARPROT   ( m_axi_gmem1_1_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_1_ARPROT
        .m_axi_gmem1_1_ARQOS    ( m_axi_gmem1_1_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_1_ARQOS
        .m_axi_gmem1_1_ARVALID  ( m_axi_gmem1_1_ARVALID  ) , // output wire m_axi_gmem1_1_ARVALID
        .m_axi_gmem1_1_ARREADY  ( m_axi_gmem1_1_ARREADY  ) , // input wire m_axi_gmem1_1_ARREADY
        .m_axi_gmem1_1_RDATA    ( m_axi_gmem1_1_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_1_RDATA
        .m_axi_gmem1_1_RRESP    ( m_axi_gmem1_1_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_1_RRESP
        .m_axi_gmem1_1_RLAST    ( m_axi_gmem1_1_RLAST    ) , // input wire m_axi_gmem1_1_RLAST
        .m_axi_gmem1_1_RVALID   ( m_axi_gmem1_1_RVALID   ) , // input wire m_axi_gmem1_1_RVALID
        .m_axi_gmem1_1_RREADY   ( m_axi_gmem1_1_RREADY   ) , // output wire m_axi_gmem1_1_RREADY
        .m_axi_gmem1_2_AWADDR   ( m_axi_gmem1_2_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_2_AWADDR
        .m_axi_gmem1_2_AWLEN    ( m_axi_gmem1_2_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_2_AWLEN
        .m_axi_gmem1_2_AWSIZE   ( m_axi_gmem1_2_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_2_AWSIZE
        .m_axi_gmem1_2_AWBURST  ( m_axi_gmem1_2_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_2_AWBURST
        .m_axi_gmem1_2_AWLOCK   ( m_axi_gmem1_2_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_2_AWLOCK
        .m_axi_gmem1_2_AWREGION ( m_axi_gmem1_2_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_2_AWREGION
        .m_axi_gmem1_2_AWCACHE  ( m_axi_gmem1_2_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_2_AWCACHE
        .m_axi_gmem1_2_AWPROT   ( m_axi_gmem1_2_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_2_AWPROT
        .m_axi_gmem1_2_AWQOS    ( m_axi_gmem1_2_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_2_AWQOS
        .m_axi_gmem1_2_AWVALID  ( m_axi_gmem1_2_AWVALID  ) , // output wire m_axi_gmem1_2_AWVALID
        .m_axi_gmem1_2_AWREADY  ( m_axi_gmem1_2_AWREADY  ) , // input wire m_axi_gmem1_2_AWREADY
        .m_axi_gmem1_2_WDATA    ( m_axi_gmem1_2_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_2_WDATA
        .m_axi_gmem1_2_WSTRB    ( m_axi_gmem1_2_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_2_WSTRB
        .m_axi_gmem1_2_WLAST    ( m_axi_gmem1_2_WLAST    ) , // output wire m_axi_gmem1_2_WLAST
        .m_axi_gmem1_2_WVALID   ( m_axi_gmem1_2_WVALID   ) , // output wire m_axi_gmem1_2_WVALID
        .m_axi_gmem1_2_WREADY   ( m_axi_gmem1_2_WREADY   ) , // input wire m_axi_gmem1_2_WREADY
        .m_axi_gmem1_2_BRESP    ( m_axi_gmem1_2_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_2_BRESP
        .m_axi_gmem1_2_BVALID   ( m_axi_gmem1_2_BVALID   ) , // input wire m_axi_gmem1_2_BVALID
        .m_axi_gmem1_2_BREADY   ( m_axi_gmem1_2_BREADY   ) , // output wire m_axi_gmem1_2_BREADY
        .m_axi_gmem1_2_ARADDR   ( m_axi_gmem1_2_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_2_ARADDR
        .m_axi_gmem1_2_ARLEN    ( m_axi_gmem1_2_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_2_ARLEN
        .m_axi_gmem1_2_ARSIZE   ( m_axi_gmem1_2_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_2_ARSIZE
        .m_axi_gmem1_2_ARBURST  ( m_axi_gmem1_2_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_2_ARBURST
        .m_axi_gmem1_2_ARLOCK   ( m_axi_gmem1_2_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_2_ARLOCK
        .m_axi_gmem1_2_ARREGION ( m_axi_gmem1_2_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_2_ARREGION
        .m_axi_gmem1_2_ARCACHE  ( m_axi_gmem1_2_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_2_ARCACHE
        .m_axi_gmem1_2_ARPROT   ( m_axi_gmem1_2_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_2_ARPROT
        .m_axi_gmem1_2_ARQOS    ( m_axi_gmem1_2_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_2_ARQOS
        .m_axi_gmem1_2_ARVALID  ( m_axi_gmem1_2_ARVALID  ) , // output wire m_axi_gmem1_2_ARVALID
        .m_axi_gmem1_2_ARREADY  ( m_axi_gmem1_2_ARREADY  ) , // input wire m_axi_gmem1_2_ARREADY
        .m_axi_gmem1_2_RDATA    ( m_axi_gmem1_2_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_2_RDATA
        .m_axi_gmem1_2_RRESP    ( m_axi_gmem1_2_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_2_RRESP
        .m_axi_gmem1_2_RLAST    ( m_axi_gmem1_2_RLAST    ) , // input wire m_axi_gmem1_2_RLAST
        .m_axi_gmem1_2_RVALID   ( m_axi_gmem1_2_RVALID   ) , // input wire m_axi_gmem1_2_RVALID
        .m_axi_gmem1_2_RREADY   ( m_axi_gmem1_2_RREADY   ) , // output wire m_axi_gmem1_2_RREADY
        .m_axi_gmem1_3_AWADDR   ( m_axi_gmem1_3_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_3_AWADDR
        .m_axi_gmem1_3_AWLEN    ( m_axi_gmem1_3_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_3_AWLEN
        .m_axi_gmem1_3_AWSIZE   ( m_axi_gmem1_3_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_3_AWSIZE
        .m_axi_gmem1_3_AWBURST  ( m_axi_gmem1_3_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_3_AWBURST
        .m_axi_gmem1_3_AWLOCK   ( m_axi_gmem1_3_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_3_AWLOCK
        .m_axi_gmem1_3_AWREGION ( m_axi_gmem1_3_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_3_AWREGION
        .m_axi_gmem1_3_AWCACHE  ( m_axi_gmem1_3_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_3_AWCACHE
        .m_axi_gmem1_3_AWPROT   ( m_axi_gmem1_3_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_3_AWPROT
        .m_axi_gmem1_3_AWQOS    ( m_axi_gmem1_3_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_3_AWQOS
        .m_axi_gmem1_3_AWVALID  ( m_axi_gmem1_3_AWVALID  ) , // output wire m_axi_gmem1_3_AWVALID
        .m_axi_gmem1_3_AWREADY  ( m_axi_gmem1_3_AWREADY  ) , // input wire m_axi_gmem1_3_AWREADY
        .m_axi_gmem1_3_WDATA    ( m_axi_gmem1_3_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_3_WDATA
        .m_axi_gmem1_3_WSTRB    ( m_axi_gmem1_3_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_3_WSTRB
        .m_axi_gmem1_3_WLAST    ( m_axi_gmem1_3_WLAST    ) , // output wire m_axi_gmem1_3_WLAST
        .m_axi_gmem1_3_WVALID   ( m_axi_gmem1_3_WVALID   ) , // output wire m_axi_gmem1_3_WVALID
        .m_axi_gmem1_3_WREADY   ( m_axi_gmem1_3_WREADY   ) , // input wire m_axi_gmem1_3_WREADY
        .m_axi_gmem1_3_BRESP    ( m_axi_gmem1_3_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_3_BRESP
        .m_axi_gmem1_3_BVALID   ( m_axi_gmem1_3_BVALID   ) , // input wire m_axi_gmem1_3_BVALID
        .m_axi_gmem1_3_BREADY   ( m_axi_gmem1_3_BREADY   ) , // output wire m_axi_gmem1_3_BREADY
        .m_axi_gmem1_3_ARADDR   ( m_axi_gmem1_3_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_3_ARADDR
        .m_axi_gmem1_3_ARLEN    ( m_axi_gmem1_3_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_3_ARLEN
        .m_axi_gmem1_3_ARSIZE   ( m_axi_gmem1_3_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_3_ARSIZE
        .m_axi_gmem1_3_ARBURST  ( m_axi_gmem1_3_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_3_ARBURST
        .m_axi_gmem1_3_ARLOCK   ( m_axi_gmem1_3_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_3_ARLOCK
        .m_axi_gmem1_3_ARREGION ( m_axi_gmem1_3_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_3_ARREGION
        .m_axi_gmem1_3_ARCACHE  ( m_axi_gmem1_3_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_3_ARCACHE
        .m_axi_gmem1_3_ARPROT   ( m_axi_gmem1_3_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_3_ARPROT
        .m_axi_gmem1_3_ARQOS    ( m_axi_gmem1_3_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_3_ARQOS
        .m_axi_gmem1_3_ARVALID  ( m_axi_gmem1_3_ARVALID  ) , // output wire m_axi_gmem1_3_ARVALID
        .m_axi_gmem1_3_ARREADY  ( m_axi_gmem1_3_ARREADY  ) , // input wire m_axi_gmem1_3_ARREADY
        .m_axi_gmem1_3_RDATA    ( m_axi_gmem1_3_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_3_RDATA
        .m_axi_gmem1_3_RRESP    ( m_axi_gmem1_3_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_3_RRESP
        .m_axi_gmem1_3_RLAST    ( m_axi_gmem1_3_RLAST    ) , // input wire m_axi_gmem1_3_RLAST
        .m_axi_gmem1_3_RVALID   ( m_axi_gmem1_3_RVALID   ) , // input wire m_axi_gmem1_3_RVALID
        .m_axi_gmem1_3_RREADY   ( m_axi_gmem1_3_RREADY   ) , // output wire m_axi_gmem1_3_RREADY
        .m_axi_gmem1_4_AWADDR   ( m_axi_gmem1_4_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_4_AWADDR
        .m_axi_gmem1_4_AWLEN    ( m_axi_gmem1_4_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_4_AWLEN
        .m_axi_gmem1_4_AWSIZE   ( m_axi_gmem1_4_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_4_AWSIZE
        .m_axi_gmem1_4_AWBURST  ( m_axi_gmem1_4_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_4_AWBURST
        .m_axi_gmem1_4_AWLOCK   ( m_axi_gmem1_4_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_4_AWLOCK
        .m_axi_gmem1_4_AWREGION ( m_axi_gmem1_4_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_4_AWREGION
        .m_axi_gmem1_4_AWCACHE  ( m_axi_gmem1_4_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_4_AWCACHE
        .m_axi_gmem1_4_AWPROT   ( m_axi_gmem1_4_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_4_AWPROT
        .m_axi_gmem1_4_AWQOS    ( m_axi_gmem1_4_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_4_AWQOS
        .m_axi_gmem1_4_AWVALID  ( m_axi_gmem1_4_AWVALID  ) , // output wire m_axi_gmem1_4_AWVALID
        .m_axi_gmem1_4_AWREADY  ( m_axi_gmem1_4_AWREADY  ) , // input wire m_axi_gmem1_4_AWREADY
        .m_axi_gmem1_4_WDATA    ( m_axi_gmem1_4_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_4_WDATA
        .m_axi_gmem1_4_WSTRB    ( m_axi_gmem1_4_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_4_WSTRB
        .m_axi_gmem1_4_WLAST    ( m_axi_gmem1_4_WLAST    ) , // output wire m_axi_gmem1_4_WLAST
        .m_axi_gmem1_4_WVALID   ( m_axi_gmem1_4_WVALID   ) , // output wire m_axi_gmem1_4_WVALID
        .m_axi_gmem1_4_WREADY   ( m_axi_gmem1_4_WREADY   ) , // input wire m_axi_gmem1_4_WREADY
        .m_axi_gmem1_4_BRESP    ( m_axi_gmem1_4_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_4_BRESP
        .m_axi_gmem1_4_BVALID   ( m_axi_gmem1_4_BVALID   ) , // input wire m_axi_gmem1_4_BVALID
        .m_axi_gmem1_4_BREADY   ( m_axi_gmem1_4_BREADY   ) , // output wire m_axi_gmem1_4_BREADY
        .m_axi_gmem1_4_ARADDR   ( m_axi_gmem1_4_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_4_ARADDR
        .m_axi_gmem1_4_ARLEN    ( m_axi_gmem1_4_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_4_ARLEN
        .m_axi_gmem1_4_ARSIZE   ( m_axi_gmem1_4_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_4_ARSIZE
        .m_axi_gmem1_4_ARBURST  ( m_axi_gmem1_4_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_4_ARBURST
        .m_axi_gmem1_4_ARLOCK   ( m_axi_gmem1_4_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_4_ARLOCK
        .m_axi_gmem1_4_ARREGION ( m_axi_gmem1_4_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_4_ARREGION
        .m_axi_gmem1_4_ARCACHE  ( m_axi_gmem1_4_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_4_ARCACHE
        .m_axi_gmem1_4_ARPROT   ( m_axi_gmem1_4_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_4_ARPROT
        .m_axi_gmem1_4_ARQOS    ( m_axi_gmem1_4_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_4_ARQOS
        .m_axi_gmem1_4_ARVALID  ( m_axi_gmem1_4_ARVALID  ) , // output wire m_axi_gmem1_4_ARVALID
        .m_axi_gmem1_4_ARREADY  ( m_axi_gmem1_4_ARREADY  ) , // input wire m_axi_gmem1_4_ARREADY
        .m_axi_gmem1_4_RDATA    ( m_axi_gmem1_4_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_4_RDATA
        .m_axi_gmem1_4_RRESP    ( m_axi_gmem1_4_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_4_RRESP
        .m_axi_gmem1_4_RLAST    ( m_axi_gmem1_4_RLAST    ) , // input wire m_axi_gmem1_4_RLAST
        .m_axi_gmem1_4_RVALID   ( m_axi_gmem1_4_RVALID   ) , // input wire m_axi_gmem1_4_RVALID
        .m_axi_gmem1_4_RREADY   ( m_axi_gmem1_4_RREADY   ) , // output wire m_axi_gmem1_4_RREADY
        .m_axi_gmem1_5_AWADDR   ( m_axi_gmem1_5_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_5_AWADDR
        .m_axi_gmem1_5_AWLEN    ( m_axi_gmem1_5_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_5_AWLEN
        .m_axi_gmem1_5_AWSIZE   ( m_axi_gmem1_5_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_5_AWSIZE
        .m_axi_gmem1_5_AWBURST  ( m_axi_gmem1_5_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_5_AWBURST
        .m_axi_gmem1_5_AWLOCK   ( m_axi_gmem1_5_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_5_AWLOCK
        .m_axi_gmem1_5_AWREGION ( m_axi_gmem1_5_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_5_AWREGION
        .m_axi_gmem1_5_AWCACHE  ( m_axi_gmem1_5_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_5_AWCACHE
        .m_axi_gmem1_5_AWPROT   ( m_axi_gmem1_5_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_5_AWPROT
        .m_axi_gmem1_5_AWQOS    ( m_axi_gmem1_5_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_5_AWQOS
        .m_axi_gmem1_5_AWVALID  ( m_axi_gmem1_5_AWVALID  ) , // output wire m_axi_gmem1_5_AWVALID
        .m_axi_gmem1_5_AWREADY  ( m_axi_gmem1_5_AWREADY  ) , // input wire m_axi_gmem1_5_AWREADY
        .m_axi_gmem1_5_WDATA    ( m_axi_gmem1_5_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_5_WDATA
        .m_axi_gmem1_5_WSTRB    ( m_axi_gmem1_5_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_5_WSTRB
        .m_axi_gmem1_5_WLAST    ( m_axi_gmem1_5_WLAST    ) , // output wire m_axi_gmem1_5_WLAST
        .m_axi_gmem1_5_WVALID   ( m_axi_gmem1_5_WVALID   ) , // output wire m_axi_gmem1_5_WVALID
        .m_axi_gmem1_5_WREADY   ( m_axi_gmem1_5_WREADY   ) , // input wire m_axi_gmem1_5_WREADY
        .m_axi_gmem1_5_BRESP    ( m_axi_gmem1_5_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_5_BRESP
        .m_axi_gmem1_5_BVALID   ( m_axi_gmem1_5_BVALID   ) , // input wire m_axi_gmem1_5_BVALID
        .m_axi_gmem1_5_BREADY   ( m_axi_gmem1_5_BREADY   ) , // output wire m_axi_gmem1_5_BREADY
        .m_axi_gmem1_5_ARADDR   ( m_axi_gmem1_5_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_5_ARADDR
        .m_axi_gmem1_5_ARLEN    ( m_axi_gmem1_5_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_5_ARLEN
        .m_axi_gmem1_5_ARSIZE   ( m_axi_gmem1_5_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_5_ARSIZE
        .m_axi_gmem1_5_ARBURST  ( m_axi_gmem1_5_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_5_ARBURST
        .m_axi_gmem1_5_ARLOCK   ( m_axi_gmem1_5_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_5_ARLOCK
        .m_axi_gmem1_5_ARREGION ( m_axi_gmem1_5_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_5_ARREGION
        .m_axi_gmem1_5_ARCACHE  ( m_axi_gmem1_5_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_5_ARCACHE
        .m_axi_gmem1_5_ARPROT   ( m_axi_gmem1_5_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_5_ARPROT
        .m_axi_gmem1_5_ARQOS    ( m_axi_gmem1_5_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_5_ARQOS
        .m_axi_gmem1_5_ARVALID  ( m_axi_gmem1_5_ARVALID  ) , // output wire m_axi_gmem1_5_ARVALID
        .m_axi_gmem1_5_ARREADY  ( m_axi_gmem1_5_ARREADY  ) , // input wire m_axi_gmem1_5_ARREADY
        .m_axi_gmem1_5_RDATA    ( m_axi_gmem1_5_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_5_RDATA
        .m_axi_gmem1_5_RRESP    ( m_axi_gmem1_5_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_5_RRESP
        .m_axi_gmem1_5_RLAST    ( m_axi_gmem1_5_RLAST    ) , // input wire m_axi_gmem1_5_RLAST
        .m_axi_gmem1_5_RVALID   ( m_axi_gmem1_5_RVALID   ) , // input wire m_axi_gmem1_5_RVALID
        .m_axi_gmem1_5_RREADY   ( m_axi_gmem1_5_RREADY   ) , // output wire m_axi_gmem1_5_RREADY
        .m_axi_gmem1_6_AWADDR   ( m_axi_gmem1_6_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_6_AWADDR
        .m_axi_gmem1_6_AWLEN    ( m_axi_gmem1_6_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_6_AWLEN
        .m_axi_gmem1_6_AWSIZE   ( m_axi_gmem1_6_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_6_AWSIZE
        .m_axi_gmem1_6_AWBURST  ( m_axi_gmem1_6_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_6_AWBURST
        .m_axi_gmem1_6_AWLOCK   ( m_axi_gmem1_6_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_6_AWLOCK
        .m_axi_gmem1_6_AWREGION ( m_axi_gmem1_6_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_6_AWREGION
        .m_axi_gmem1_6_AWCACHE  ( m_axi_gmem1_6_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_6_AWCACHE
        .m_axi_gmem1_6_AWPROT   ( m_axi_gmem1_6_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_6_AWPROT
        .m_axi_gmem1_6_AWQOS    ( m_axi_gmem1_6_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_6_AWQOS
        .m_axi_gmem1_6_AWVALID  ( m_axi_gmem1_6_AWVALID  ) , // output wire m_axi_gmem1_6_AWVALID
        .m_axi_gmem1_6_AWREADY  ( m_axi_gmem1_6_AWREADY  ) , // input wire m_axi_gmem1_6_AWREADY
        .m_axi_gmem1_6_WDATA    ( m_axi_gmem1_6_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_6_WDATA
        .m_axi_gmem1_6_WSTRB    ( m_axi_gmem1_6_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_6_WSTRB
        .m_axi_gmem1_6_WLAST    ( m_axi_gmem1_6_WLAST    ) , // output wire m_axi_gmem1_6_WLAST
        .m_axi_gmem1_6_WVALID   ( m_axi_gmem1_6_WVALID   ) , // output wire m_axi_gmem1_6_WVALID
        .m_axi_gmem1_6_WREADY   ( m_axi_gmem1_6_WREADY   ) , // input wire m_axi_gmem1_6_WREADY
        .m_axi_gmem1_6_BRESP    ( m_axi_gmem1_6_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_6_BRESP
        .m_axi_gmem1_6_BVALID   ( m_axi_gmem1_6_BVALID   ) , // input wire m_axi_gmem1_6_BVALID
        .m_axi_gmem1_6_BREADY   ( m_axi_gmem1_6_BREADY   ) , // output wire m_axi_gmem1_6_BREADY
        .m_axi_gmem1_6_ARADDR   ( m_axi_gmem1_6_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_6_ARADDR
        .m_axi_gmem1_6_ARLEN    ( m_axi_gmem1_6_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_6_ARLEN
        .m_axi_gmem1_6_ARSIZE   ( m_axi_gmem1_6_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_6_ARSIZE
        .m_axi_gmem1_6_ARBURST  ( m_axi_gmem1_6_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_6_ARBURST
        .m_axi_gmem1_6_ARLOCK   ( m_axi_gmem1_6_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_6_ARLOCK
        .m_axi_gmem1_6_ARREGION ( m_axi_gmem1_6_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_6_ARREGION
        .m_axi_gmem1_6_ARCACHE  ( m_axi_gmem1_6_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_6_ARCACHE
        .m_axi_gmem1_6_ARPROT   ( m_axi_gmem1_6_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_6_ARPROT
        .m_axi_gmem1_6_ARQOS    ( m_axi_gmem1_6_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_6_ARQOS
        .m_axi_gmem1_6_ARVALID  ( m_axi_gmem1_6_ARVALID  ) , // output wire m_axi_gmem1_6_ARVALID
        .m_axi_gmem1_6_ARREADY  ( m_axi_gmem1_6_ARREADY  ) , // input wire m_axi_gmem1_6_ARREADY
        .m_axi_gmem1_6_RDATA    ( m_axi_gmem1_6_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_6_RDATA
        .m_axi_gmem1_6_RRESP    ( m_axi_gmem1_6_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_6_RRESP
        .m_axi_gmem1_6_RLAST    ( m_axi_gmem1_6_RLAST    ) , // input wire m_axi_gmem1_6_RLAST
        .m_axi_gmem1_6_RVALID   ( m_axi_gmem1_6_RVALID   ) , // input wire m_axi_gmem1_6_RVALID
        .m_axi_gmem1_6_RREADY   ( m_axi_gmem1_6_RREADY   ) , // output wire m_axi_gmem1_6_RREADY
        .m_axi_gmem1_7_AWADDR   ( m_axi_gmem1_7_AWADDR   ) , // output wire [63 : 0] m_axi_gmem1_7_AWADDR
        .m_axi_gmem1_7_AWLEN    ( m_axi_gmem1_7_AWLEN    ) , // output wire [7 : 0] m_axi_gmem1_7_AWLEN
        .m_axi_gmem1_7_AWSIZE   ( m_axi_gmem1_7_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem1_7_AWSIZE
        .m_axi_gmem1_7_AWBURST  ( m_axi_gmem1_7_AWBURST  ) , // output wire [1 : 0] m_axi_gmem1_7_AWBURST
        .m_axi_gmem1_7_AWLOCK   ( m_axi_gmem1_7_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem1_7_AWLOCK
        .m_axi_gmem1_7_AWREGION ( m_axi_gmem1_7_AWREGION ) , // output wire [3 : 0] m_axi_gmem1_7_AWREGION
        .m_axi_gmem1_7_AWCACHE  ( m_axi_gmem1_7_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem1_7_AWCACHE
        .m_axi_gmem1_7_AWPROT   ( m_axi_gmem1_7_AWPROT   ) , // output wire [2 : 0] m_axi_gmem1_7_AWPROT
        .m_axi_gmem1_7_AWQOS    ( m_axi_gmem1_7_AWQOS    ) , // output wire [3 : 0] m_axi_gmem1_7_AWQOS
        .m_axi_gmem1_7_AWVALID  ( m_axi_gmem1_7_AWVALID  ) , // output wire m_axi_gmem1_7_AWVALID
        .m_axi_gmem1_7_AWREADY  ( m_axi_gmem1_7_AWREADY  ) , // input wire m_axi_gmem1_7_AWREADY
        .m_axi_gmem1_7_WDATA    ( m_axi_gmem1_7_WDATA    ) , // output wire [63 : 0] m_axi_gmem1_7_WDATA
        .m_axi_gmem1_7_WSTRB    ( m_axi_gmem1_7_WSTRB    ) , // output wire [7 : 0] m_axi_gmem1_7_WSTRB
        .m_axi_gmem1_7_WLAST    ( m_axi_gmem1_7_WLAST    ) , // output wire m_axi_gmem1_7_WLAST
        .m_axi_gmem1_7_WVALID   ( m_axi_gmem1_7_WVALID   ) , // output wire m_axi_gmem1_7_WVALID
        .m_axi_gmem1_7_WREADY   ( m_axi_gmem1_7_WREADY   ) , // input wire m_axi_gmem1_7_WREADY
        .m_axi_gmem1_7_BRESP    ( m_axi_gmem1_7_BRESP    ) , // input wire [1 : 0] m_axi_gmem1_7_BRESP
        .m_axi_gmem1_7_BVALID   ( m_axi_gmem1_7_BVALID   ) , // input wire m_axi_gmem1_7_BVALID
        .m_axi_gmem1_7_BREADY   ( m_axi_gmem1_7_BREADY   ) , // output wire m_axi_gmem1_7_BREADY
        .m_axi_gmem1_7_ARADDR   ( m_axi_gmem1_7_ARADDR   ) , // output wire [63 : 0] m_axi_gmem1_7_ARADDR
        .m_axi_gmem1_7_ARLEN    ( m_axi_gmem1_7_ARLEN    ) , // output wire [7 : 0] m_axi_gmem1_7_ARLEN
        .m_axi_gmem1_7_ARSIZE   ( m_axi_gmem1_7_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem1_7_ARSIZE
        .m_axi_gmem1_7_ARBURST  ( m_axi_gmem1_7_ARBURST  ) , // output wire [1 : 0] m_axi_gmem1_7_ARBURST
        .m_axi_gmem1_7_ARLOCK   ( m_axi_gmem1_7_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem1_7_ARLOCK
        .m_axi_gmem1_7_ARREGION ( m_axi_gmem1_7_ARREGION ) , // output wire [3 : 0] m_axi_gmem1_7_ARREGION
        .m_axi_gmem1_7_ARCACHE  ( m_axi_gmem1_7_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem1_7_ARCACHE
        .m_axi_gmem1_7_ARPROT   ( m_axi_gmem1_7_ARPROT   ) , // output wire [2 : 0] m_axi_gmem1_7_ARPROT
        .m_axi_gmem1_7_ARQOS    ( m_axi_gmem1_7_ARQOS    ) , // output wire [3 : 0] m_axi_gmem1_7_ARQOS
        .m_axi_gmem1_7_ARVALID  ( m_axi_gmem1_7_ARVALID  ) , // output wire m_axi_gmem1_7_ARVALID
        .m_axi_gmem1_7_ARREADY  ( m_axi_gmem1_7_ARREADY  ) , // input wire m_axi_gmem1_7_ARREADY
        .m_axi_gmem1_7_RDATA    ( m_axi_gmem1_7_RDATA    ) , // input wire [63 : 0] m_axi_gmem1_7_RDATA
        .m_axi_gmem1_7_RRESP    ( m_axi_gmem1_7_RRESP    ) , // input wire [1 : 0] m_axi_gmem1_7_RRESP
        .m_axi_gmem1_7_RLAST    ( m_axi_gmem1_7_RLAST    ) , // input wire m_axi_gmem1_7_RLAST
        .m_axi_gmem1_7_RVALID   ( m_axi_gmem1_7_RVALID   ) , // input wire m_axi_gmem1_7_RVALID
        .m_axi_gmem1_7_RREADY   ( m_axi_gmem1_7_RREADY   ) , // output wire m_axi_gmem1_7_RREADY
        .m_axi_gmem2_0_AWADDR   ( m_axi_gmem2_0_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_0_AWADDR
        .m_axi_gmem2_0_AWLEN    ( m_axi_gmem2_0_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_0_AWLEN
        .m_axi_gmem2_0_AWSIZE   ( m_axi_gmem2_0_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_0_AWSIZE
        .m_axi_gmem2_0_AWBURST  ( m_axi_gmem2_0_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_0_AWBURST
        .m_axi_gmem2_0_AWLOCK   ( m_axi_gmem2_0_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_0_AWLOCK
        .m_axi_gmem2_0_AWREGION ( m_axi_gmem2_0_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_0_AWREGION
        .m_axi_gmem2_0_AWCACHE  ( m_axi_gmem2_0_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_0_AWCACHE
        .m_axi_gmem2_0_AWPROT   ( m_axi_gmem2_0_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_0_AWPROT
        .m_axi_gmem2_0_AWQOS    ( m_axi_gmem2_0_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_0_AWQOS
        .m_axi_gmem2_0_AWVALID  ( m_axi_gmem2_0_AWVALID  ) , // output wire m_axi_gmem2_0_AWVALID
        .m_axi_gmem2_0_AWREADY  ( m_axi_gmem2_0_AWREADY  ) , // input wire m_axi_gmem2_0_AWREADY
        .m_axi_gmem2_0_WDATA    ( m_axi_gmem2_0_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_0_WDATA
        .m_axi_gmem2_0_WSTRB    ( m_axi_gmem2_0_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_0_WSTRB
        .m_axi_gmem2_0_WLAST    ( m_axi_gmem2_0_WLAST    ) , // output wire m_axi_gmem2_0_WLAST
        .m_axi_gmem2_0_WVALID   ( m_axi_gmem2_0_WVALID   ) , // output wire m_axi_gmem2_0_WVALID
        .m_axi_gmem2_0_WREADY   ( m_axi_gmem2_0_WREADY   ) , // input wire m_axi_gmem2_0_WREADY
        .m_axi_gmem2_0_BRESP    ( m_axi_gmem2_0_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_0_BRESP
        .m_axi_gmem2_0_BVALID   ( m_axi_gmem2_0_BVALID   ) , // input wire m_axi_gmem2_0_BVALID
        .m_axi_gmem2_0_BREADY   ( m_axi_gmem2_0_BREADY   ) , // output wire m_axi_gmem2_0_BREADY
        .m_axi_gmem2_0_ARADDR   ( m_axi_gmem2_0_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_0_ARADDR
        .m_axi_gmem2_0_ARLEN    ( m_axi_gmem2_0_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_0_ARLEN
        .m_axi_gmem2_0_ARSIZE   ( m_axi_gmem2_0_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_0_ARSIZE
        .m_axi_gmem2_0_ARBURST  ( m_axi_gmem2_0_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_0_ARBURST
        .m_axi_gmem2_0_ARLOCK   ( m_axi_gmem2_0_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_0_ARLOCK
        .m_axi_gmem2_0_ARREGION ( m_axi_gmem2_0_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_0_ARREGION
        .m_axi_gmem2_0_ARCACHE  ( m_axi_gmem2_0_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_0_ARCACHE
        .m_axi_gmem2_0_ARPROT   ( m_axi_gmem2_0_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_0_ARPROT
        .m_axi_gmem2_0_ARQOS    ( m_axi_gmem2_0_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_0_ARQOS
        .m_axi_gmem2_0_ARVALID  ( m_axi_gmem2_0_ARVALID  ) , // output wire m_axi_gmem2_0_ARVALID
        .m_axi_gmem2_0_ARREADY  ( m_axi_gmem2_0_ARREADY  ) , // input wire m_axi_gmem2_0_ARREADY
        .m_axi_gmem2_0_RDATA    ( m_axi_gmem2_0_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_0_RDATA
        .m_axi_gmem2_0_RRESP    ( m_axi_gmem2_0_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_0_RRESP
        .m_axi_gmem2_0_RLAST    ( m_axi_gmem2_0_RLAST    ) , // input wire m_axi_gmem2_0_RLAST
        .m_axi_gmem2_0_RVALID   ( m_axi_gmem2_0_RVALID   ) , // input wire m_axi_gmem2_0_RVALID
        .m_axi_gmem2_0_RREADY   ( m_axi_gmem2_0_RREADY   ) , // output wire m_axi_gmem2_0_RREADY
        .m_axi_gmem2_1_AWADDR   ( m_axi_gmem2_1_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_1_AWADDR
        .m_axi_gmem2_1_AWLEN    ( m_axi_gmem2_1_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_1_AWLEN
        .m_axi_gmem2_1_AWSIZE   ( m_axi_gmem2_1_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_1_AWSIZE
        .m_axi_gmem2_1_AWBURST  ( m_axi_gmem2_1_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_1_AWBURST
        .m_axi_gmem2_1_AWLOCK   ( m_axi_gmem2_1_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_1_AWLOCK
        .m_axi_gmem2_1_AWREGION ( m_axi_gmem2_1_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_1_AWREGION
        .m_axi_gmem2_1_AWCACHE  ( m_axi_gmem2_1_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_1_AWCACHE
        .m_axi_gmem2_1_AWPROT   ( m_axi_gmem2_1_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_1_AWPROT
        .m_axi_gmem2_1_AWQOS    ( m_axi_gmem2_1_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_1_AWQOS
        .m_axi_gmem2_1_AWVALID  ( m_axi_gmem2_1_AWVALID  ) , // output wire m_axi_gmem2_1_AWVALID
        .m_axi_gmem2_1_AWREADY  ( m_axi_gmem2_1_AWREADY  ) , // input wire m_axi_gmem2_1_AWREADY
        .m_axi_gmem2_1_WDATA    ( m_axi_gmem2_1_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_1_WDATA
        .m_axi_gmem2_1_WSTRB    ( m_axi_gmem2_1_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_1_WSTRB
        .m_axi_gmem2_1_WLAST    ( m_axi_gmem2_1_WLAST    ) , // output wire m_axi_gmem2_1_WLAST
        .m_axi_gmem2_1_WVALID   ( m_axi_gmem2_1_WVALID   ) , // output wire m_axi_gmem2_1_WVALID
        .m_axi_gmem2_1_WREADY   ( m_axi_gmem2_1_WREADY   ) , // input wire m_axi_gmem2_1_WREADY
        .m_axi_gmem2_1_BRESP    ( m_axi_gmem2_1_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_1_BRESP
        .m_axi_gmem2_1_BVALID   ( m_axi_gmem2_1_BVALID   ) , // input wire m_axi_gmem2_1_BVALID
        .m_axi_gmem2_1_BREADY   ( m_axi_gmem2_1_BREADY   ) , // output wire m_axi_gmem2_1_BREADY
        .m_axi_gmem2_1_ARADDR   ( m_axi_gmem2_1_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_1_ARADDR
        .m_axi_gmem2_1_ARLEN    ( m_axi_gmem2_1_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_1_ARLEN
        .m_axi_gmem2_1_ARSIZE   ( m_axi_gmem2_1_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_1_ARSIZE
        .m_axi_gmem2_1_ARBURST  ( m_axi_gmem2_1_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_1_ARBURST
        .m_axi_gmem2_1_ARLOCK   ( m_axi_gmem2_1_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_1_ARLOCK
        .m_axi_gmem2_1_ARREGION ( m_axi_gmem2_1_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_1_ARREGION
        .m_axi_gmem2_1_ARCACHE  ( m_axi_gmem2_1_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_1_ARCACHE
        .m_axi_gmem2_1_ARPROT   ( m_axi_gmem2_1_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_1_ARPROT
        .m_axi_gmem2_1_ARQOS    ( m_axi_gmem2_1_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_1_ARQOS
        .m_axi_gmem2_1_ARVALID  ( m_axi_gmem2_1_ARVALID  ) , // output wire m_axi_gmem2_1_ARVALID
        .m_axi_gmem2_1_ARREADY  ( m_axi_gmem2_1_ARREADY  ) , // input wire m_axi_gmem2_1_ARREADY
        .m_axi_gmem2_1_RDATA    ( m_axi_gmem2_1_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_1_RDATA
        .m_axi_gmem2_1_RRESP    ( m_axi_gmem2_1_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_1_RRESP
        .m_axi_gmem2_1_RLAST    ( m_axi_gmem2_1_RLAST    ) , // input wire m_axi_gmem2_1_RLAST
        .m_axi_gmem2_1_RVALID   ( m_axi_gmem2_1_RVALID   ) , // input wire m_axi_gmem2_1_RVALID
        .m_axi_gmem2_1_RREADY   ( m_axi_gmem2_1_RREADY   ) , // output wire m_axi_gmem2_1_RREADY
        .m_axi_gmem2_2_AWADDR   ( m_axi_gmem2_2_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_2_AWADDR
        .m_axi_gmem2_2_AWLEN    ( m_axi_gmem2_2_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_2_AWLEN
        .m_axi_gmem2_2_AWSIZE   ( m_axi_gmem2_2_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_2_AWSIZE
        .m_axi_gmem2_2_AWBURST  ( m_axi_gmem2_2_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_2_AWBURST
        .m_axi_gmem2_2_AWLOCK   ( m_axi_gmem2_2_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_2_AWLOCK
        .m_axi_gmem2_2_AWREGION ( m_axi_gmem2_2_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_2_AWREGION
        .m_axi_gmem2_2_AWCACHE  ( m_axi_gmem2_2_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_2_AWCACHE
        .m_axi_gmem2_2_AWPROT   ( m_axi_gmem2_2_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_2_AWPROT
        .m_axi_gmem2_2_AWQOS    ( m_axi_gmem2_2_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_2_AWQOS
        .m_axi_gmem2_2_AWVALID  ( m_axi_gmem2_2_AWVALID  ) , // output wire m_axi_gmem2_2_AWVALID
        .m_axi_gmem2_2_AWREADY  ( m_axi_gmem2_2_AWREADY  ) , // input wire m_axi_gmem2_2_AWREADY
        .m_axi_gmem2_2_WDATA    ( m_axi_gmem2_2_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_2_WDATA
        .m_axi_gmem2_2_WSTRB    ( m_axi_gmem2_2_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_2_WSTRB
        .m_axi_gmem2_2_WLAST    ( m_axi_gmem2_2_WLAST    ) , // output wire m_axi_gmem2_2_WLAST
        .m_axi_gmem2_2_WVALID   ( m_axi_gmem2_2_WVALID   ) , // output wire m_axi_gmem2_2_WVALID
        .m_axi_gmem2_2_WREADY   ( m_axi_gmem2_2_WREADY   ) , // input wire m_axi_gmem2_2_WREADY
        .m_axi_gmem2_2_BRESP    ( m_axi_gmem2_2_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_2_BRESP
        .m_axi_gmem2_2_BVALID   ( m_axi_gmem2_2_BVALID   ) , // input wire m_axi_gmem2_2_BVALID
        .m_axi_gmem2_2_BREADY   ( m_axi_gmem2_2_BREADY   ) , // output wire m_axi_gmem2_2_BREADY
        .m_axi_gmem2_2_ARADDR   ( m_axi_gmem2_2_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_2_ARADDR
        .m_axi_gmem2_2_ARLEN    ( m_axi_gmem2_2_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_2_ARLEN
        .m_axi_gmem2_2_ARSIZE   ( m_axi_gmem2_2_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_2_ARSIZE
        .m_axi_gmem2_2_ARBURST  ( m_axi_gmem2_2_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_2_ARBURST
        .m_axi_gmem2_2_ARLOCK   ( m_axi_gmem2_2_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_2_ARLOCK
        .m_axi_gmem2_2_ARREGION ( m_axi_gmem2_2_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_2_ARREGION
        .m_axi_gmem2_2_ARCACHE  ( m_axi_gmem2_2_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_2_ARCACHE
        .m_axi_gmem2_2_ARPROT   ( m_axi_gmem2_2_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_2_ARPROT
        .m_axi_gmem2_2_ARQOS    ( m_axi_gmem2_2_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_2_ARQOS
        .m_axi_gmem2_2_ARVALID  ( m_axi_gmem2_2_ARVALID  ) , // output wire m_axi_gmem2_2_ARVALID
        .m_axi_gmem2_2_ARREADY  ( m_axi_gmem2_2_ARREADY  ) , // input wire m_axi_gmem2_2_ARREADY
        .m_axi_gmem2_2_RDATA    ( m_axi_gmem2_2_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_2_RDATA
        .m_axi_gmem2_2_RRESP    ( m_axi_gmem2_2_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_2_RRESP
        .m_axi_gmem2_2_RLAST    ( m_axi_gmem2_2_RLAST    ) , // input wire m_axi_gmem2_2_RLAST
        .m_axi_gmem2_2_RVALID   ( m_axi_gmem2_2_RVALID   ) , // input wire m_axi_gmem2_2_RVALID
        .m_axi_gmem2_2_RREADY   ( m_axi_gmem2_2_RREADY   ) , // output wire m_axi_gmem2_2_RREADY
        .m_axi_gmem2_3_AWADDR   ( m_axi_gmem2_3_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_3_AWADDR
        .m_axi_gmem2_3_AWLEN    ( m_axi_gmem2_3_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_3_AWLEN
        .m_axi_gmem2_3_AWSIZE   ( m_axi_gmem2_3_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_3_AWSIZE
        .m_axi_gmem2_3_AWBURST  ( m_axi_gmem2_3_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_3_AWBURST
        .m_axi_gmem2_3_AWLOCK   ( m_axi_gmem2_3_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_3_AWLOCK
        .m_axi_gmem2_3_AWREGION ( m_axi_gmem2_3_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_3_AWREGION
        .m_axi_gmem2_3_AWCACHE  ( m_axi_gmem2_3_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_3_AWCACHE
        .m_axi_gmem2_3_AWPROT   ( m_axi_gmem2_3_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_3_AWPROT
        .m_axi_gmem2_3_AWQOS    ( m_axi_gmem2_3_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_3_AWQOS
        .m_axi_gmem2_3_AWVALID  ( m_axi_gmem2_3_AWVALID  ) , // output wire m_axi_gmem2_3_AWVALID
        .m_axi_gmem2_3_AWREADY  ( m_axi_gmem2_3_AWREADY  ) , // input wire m_axi_gmem2_3_AWREADY
        .m_axi_gmem2_3_WDATA    ( m_axi_gmem2_3_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_3_WDATA
        .m_axi_gmem2_3_WSTRB    ( m_axi_gmem2_3_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_3_WSTRB
        .m_axi_gmem2_3_WLAST    ( m_axi_gmem2_3_WLAST    ) , // output wire m_axi_gmem2_3_WLAST
        .m_axi_gmem2_3_WVALID   ( m_axi_gmem2_3_WVALID   ) , // output wire m_axi_gmem2_3_WVALID
        .m_axi_gmem2_3_WREADY   ( m_axi_gmem2_3_WREADY   ) , // input wire m_axi_gmem2_3_WREADY
        .m_axi_gmem2_3_BRESP    ( m_axi_gmem2_3_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_3_BRESP
        .m_axi_gmem2_3_BVALID   ( m_axi_gmem2_3_BVALID   ) , // input wire m_axi_gmem2_3_BVALID
        .m_axi_gmem2_3_BREADY   ( m_axi_gmem2_3_BREADY   ) , // output wire m_axi_gmem2_3_BREADY
        .m_axi_gmem2_3_ARADDR   ( m_axi_gmem2_3_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_3_ARADDR
        .m_axi_gmem2_3_ARLEN    ( m_axi_gmem2_3_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_3_ARLEN
        .m_axi_gmem2_3_ARSIZE   ( m_axi_gmem2_3_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_3_ARSIZE
        .m_axi_gmem2_3_ARBURST  ( m_axi_gmem2_3_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_3_ARBURST
        .m_axi_gmem2_3_ARLOCK   ( m_axi_gmem2_3_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_3_ARLOCK
        .m_axi_gmem2_3_ARREGION ( m_axi_gmem2_3_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_3_ARREGION
        .m_axi_gmem2_3_ARCACHE  ( m_axi_gmem2_3_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_3_ARCACHE
        .m_axi_gmem2_3_ARPROT   ( m_axi_gmem2_3_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_3_ARPROT
        .m_axi_gmem2_3_ARQOS    ( m_axi_gmem2_3_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_3_ARQOS
        .m_axi_gmem2_3_ARVALID  ( m_axi_gmem2_3_ARVALID  ) , // output wire m_axi_gmem2_3_ARVALID
        .m_axi_gmem2_3_ARREADY  ( m_axi_gmem2_3_ARREADY  ) , // input wire m_axi_gmem2_3_ARREADY
        .m_axi_gmem2_3_RDATA    ( m_axi_gmem2_3_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_3_RDATA
        .m_axi_gmem2_3_RRESP    ( m_axi_gmem2_3_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_3_RRESP
        .m_axi_gmem2_3_RLAST    ( m_axi_gmem2_3_RLAST    ) , // input wire m_axi_gmem2_3_RLAST
        .m_axi_gmem2_3_RVALID   ( m_axi_gmem2_3_RVALID   ) , // input wire m_axi_gmem2_3_RVALID
        .m_axi_gmem2_3_RREADY   ( m_axi_gmem2_3_RREADY   ) , // output wire m_axi_gmem2_3_RREADY
        .m_axi_gmem2_4_AWADDR   ( m_axi_gmem2_4_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_4_AWADDR
        .m_axi_gmem2_4_AWLEN    ( m_axi_gmem2_4_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_4_AWLEN
        .m_axi_gmem2_4_AWSIZE   ( m_axi_gmem2_4_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_4_AWSIZE
        .m_axi_gmem2_4_AWBURST  ( m_axi_gmem2_4_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_4_AWBURST
        .m_axi_gmem2_4_AWLOCK   ( m_axi_gmem2_4_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_4_AWLOCK
        .m_axi_gmem2_4_AWREGION ( m_axi_gmem2_4_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_4_AWREGION
        .m_axi_gmem2_4_AWCACHE  ( m_axi_gmem2_4_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_4_AWCACHE
        .m_axi_gmem2_4_AWPROT   ( m_axi_gmem2_4_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_4_AWPROT
        .m_axi_gmem2_4_AWQOS    ( m_axi_gmem2_4_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_4_AWQOS
        .m_axi_gmem2_4_AWVALID  ( m_axi_gmem2_4_AWVALID  ) , // output wire m_axi_gmem2_4_AWVALID
        .m_axi_gmem2_4_AWREADY  ( m_axi_gmem2_4_AWREADY  ) , // input wire m_axi_gmem2_4_AWREADY
        .m_axi_gmem2_4_WDATA    ( m_axi_gmem2_4_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_4_WDATA
        .m_axi_gmem2_4_WSTRB    ( m_axi_gmem2_4_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_4_WSTRB
        .m_axi_gmem2_4_WLAST    ( m_axi_gmem2_4_WLAST    ) , // output wire m_axi_gmem2_4_WLAST
        .m_axi_gmem2_4_WVALID   ( m_axi_gmem2_4_WVALID   ) , // output wire m_axi_gmem2_4_WVALID
        .m_axi_gmem2_4_WREADY   ( m_axi_gmem2_4_WREADY   ) , // input wire m_axi_gmem2_4_WREADY
        .m_axi_gmem2_4_BRESP    ( m_axi_gmem2_4_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_4_BRESP
        .m_axi_gmem2_4_BVALID   ( m_axi_gmem2_4_BVALID   ) , // input wire m_axi_gmem2_4_BVALID
        .m_axi_gmem2_4_BREADY   ( m_axi_gmem2_4_BREADY   ) , // output wire m_axi_gmem2_4_BREADY
        .m_axi_gmem2_4_ARADDR   ( m_axi_gmem2_4_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_4_ARADDR
        .m_axi_gmem2_4_ARLEN    ( m_axi_gmem2_4_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_4_ARLEN
        .m_axi_gmem2_4_ARSIZE   ( m_axi_gmem2_4_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_4_ARSIZE
        .m_axi_gmem2_4_ARBURST  ( m_axi_gmem2_4_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_4_ARBURST
        .m_axi_gmem2_4_ARLOCK   ( m_axi_gmem2_4_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_4_ARLOCK
        .m_axi_gmem2_4_ARREGION ( m_axi_gmem2_4_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_4_ARREGION
        .m_axi_gmem2_4_ARCACHE  ( m_axi_gmem2_4_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_4_ARCACHE
        .m_axi_gmem2_4_ARPROT   ( m_axi_gmem2_4_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_4_ARPROT
        .m_axi_gmem2_4_ARQOS    ( m_axi_gmem2_4_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_4_ARQOS
        .m_axi_gmem2_4_ARVALID  ( m_axi_gmem2_4_ARVALID  ) , // output wire m_axi_gmem2_4_ARVALID
        .m_axi_gmem2_4_ARREADY  ( m_axi_gmem2_4_ARREADY  ) , // input wire m_axi_gmem2_4_ARREADY
        .m_axi_gmem2_4_RDATA    ( m_axi_gmem2_4_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_4_RDATA
        .m_axi_gmem2_4_RRESP    ( m_axi_gmem2_4_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_4_RRESP
        .m_axi_gmem2_4_RLAST    ( m_axi_gmem2_4_RLAST    ) , // input wire m_axi_gmem2_4_RLAST
        .m_axi_gmem2_4_RVALID   ( m_axi_gmem2_4_RVALID   ) , // input wire m_axi_gmem2_4_RVALID
        .m_axi_gmem2_4_RREADY   ( m_axi_gmem2_4_RREADY   ) , // output wire m_axi_gmem2_4_RREADY
        .m_axi_gmem2_5_AWADDR   ( m_axi_gmem2_5_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_5_AWADDR
        .m_axi_gmem2_5_AWLEN    ( m_axi_gmem2_5_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_5_AWLEN
        .m_axi_gmem2_5_AWSIZE   ( m_axi_gmem2_5_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_5_AWSIZE
        .m_axi_gmem2_5_AWBURST  ( m_axi_gmem2_5_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_5_AWBURST
        .m_axi_gmem2_5_AWLOCK   ( m_axi_gmem2_5_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_5_AWLOCK
        .m_axi_gmem2_5_AWREGION ( m_axi_gmem2_5_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_5_AWREGION
        .m_axi_gmem2_5_AWCACHE  ( m_axi_gmem2_5_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_5_AWCACHE
        .m_axi_gmem2_5_AWPROT   ( m_axi_gmem2_5_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_5_AWPROT
        .m_axi_gmem2_5_AWQOS    ( m_axi_gmem2_5_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_5_AWQOS
        .m_axi_gmem2_5_AWVALID  ( m_axi_gmem2_5_AWVALID  ) , // output wire m_axi_gmem2_5_AWVALID
        .m_axi_gmem2_5_AWREADY  ( m_axi_gmem2_5_AWREADY  ) , // input wire m_axi_gmem2_5_AWREADY
        .m_axi_gmem2_5_WDATA    ( m_axi_gmem2_5_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_5_WDATA
        .m_axi_gmem2_5_WSTRB    ( m_axi_gmem2_5_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_5_WSTRB
        .m_axi_gmem2_5_WLAST    ( m_axi_gmem2_5_WLAST    ) , // output wire m_axi_gmem2_5_WLAST
        .m_axi_gmem2_5_WVALID   ( m_axi_gmem2_5_WVALID   ) , // output wire m_axi_gmem2_5_WVALID
        .m_axi_gmem2_5_WREADY   ( m_axi_gmem2_5_WREADY   ) , // input wire m_axi_gmem2_5_WREADY
        .m_axi_gmem2_5_BRESP    ( m_axi_gmem2_5_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_5_BRESP
        .m_axi_gmem2_5_BVALID   ( m_axi_gmem2_5_BVALID   ) , // input wire m_axi_gmem2_5_BVALID
        .m_axi_gmem2_5_BREADY   ( m_axi_gmem2_5_BREADY   ) , // output wire m_axi_gmem2_5_BREADY
        .m_axi_gmem2_5_ARADDR   ( m_axi_gmem2_5_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_5_ARADDR
        .m_axi_gmem2_5_ARLEN    ( m_axi_gmem2_5_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_5_ARLEN
        .m_axi_gmem2_5_ARSIZE   ( m_axi_gmem2_5_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_5_ARSIZE
        .m_axi_gmem2_5_ARBURST  ( m_axi_gmem2_5_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_5_ARBURST
        .m_axi_gmem2_5_ARLOCK   ( m_axi_gmem2_5_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_5_ARLOCK
        .m_axi_gmem2_5_ARREGION ( m_axi_gmem2_5_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_5_ARREGION
        .m_axi_gmem2_5_ARCACHE  ( m_axi_gmem2_5_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_5_ARCACHE
        .m_axi_gmem2_5_ARPROT   ( m_axi_gmem2_5_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_5_ARPROT
        .m_axi_gmem2_5_ARQOS    ( m_axi_gmem2_5_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_5_ARQOS
        .m_axi_gmem2_5_ARVALID  ( m_axi_gmem2_5_ARVALID  ) , // output wire m_axi_gmem2_5_ARVALID
        .m_axi_gmem2_5_ARREADY  ( m_axi_gmem2_5_ARREADY  ) , // input wire m_axi_gmem2_5_ARREADY
        .m_axi_gmem2_5_RDATA    ( m_axi_gmem2_5_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_5_RDATA
        .m_axi_gmem2_5_RRESP    ( m_axi_gmem2_5_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_5_RRESP
        .m_axi_gmem2_5_RLAST    ( m_axi_gmem2_5_RLAST    ) , // input wire m_axi_gmem2_5_RLAST
        .m_axi_gmem2_5_RVALID   ( m_axi_gmem2_5_RVALID   ) , // input wire m_axi_gmem2_5_RVALID
        .m_axi_gmem2_5_RREADY   ( m_axi_gmem2_5_RREADY   ) , // output wire m_axi_gmem2_5_RREADY
        .m_axi_gmem2_6_AWADDR   ( m_axi_gmem2_6_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_6_AWADDR
        .m_axi_gmem2_6_AWLEN    ( m_axi_gmem2_6_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_6_AWLEN
        .m_axi_gmem2_6_AWSIZE   ( m_axi_gmem2_6_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_6_AWSIZE
        .m_axi_gmem2_6_AWBURST  ( m_axi_gmem2_6_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_6_AWBURST
        .m_axi_gmem2_6_AWLOCK   ( m_axi_gmem2_6_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_6_AWLOCK
        .m_axi_gmem2_6_AWREGION ( m_axi_gmem2_6_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_6_AWREGION
        .m_axi_gmem2_6_AWCACHE  ( m_axi_gmem2_6_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_6_AWCACHE
        .m_axi_gmem2_6_AWPROT   ( m_axi_gmem2_6_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_6_AWPROT
        .m_axi_gmem2_6_AWQOS    ( m_axi_gmem2_6_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_6_AWQOS
        .m_axi_gmem2_6_AWVALID  ( m_axi_gmem2_6_AWVALID  ) , // output wire m_axi_gmem2_6_AWVALID
        .m_axi_gmem2_6_AWREADY  ( m_axi_gmem2_6_AWREADY  ) , // input wire m_axi_gmem2_6_AWREADY
        .m_axi_gmem2_6_WDATA    ( m_axi_gmem2_6_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_6_WDATA
        .m_axi_gmem2_6_WSTRB    ( m_axi_gmem2_6_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_6_WSTRB
        .m_axi_gmem2_6_WLAST    ( m_axi_gmem2_6_WLAST    ) , // output wire m_axi_gmem2_6_WLAST
        .m_axi_gmem2_6_WVALID   ( m_axi_gmem2_6_WVALID   ) , // output wire m_axi_gmem2_6_WVALID
        .m_axi_gmem2_6_WREADY   ( m_axi_gmem2_6_WREADY   ) , // input wire m_axi_gmem2_6_WREADY
        .m_axi_gmem2_6_BRESP    ( m_axi_gmem2_6_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_6_BRESP
        .m_axi_gmem2_6_BVALID   ( m_axi_gmem2_6_BVALID   ) , // input wire m_axi_gmem2_6_BVALID
        .m_axi_gmem2_6_BREADY   ( m_axi_gmem2_6_BREADY   ) , // output wire m_axi_gmem2_6_BREADY
        .m_axi_gmem2_6_ARADDR   ( m_axi_gmem2_6_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_6_ARADDR
        .m_axi_gmem2_6_ARLEN    ( m_axi_gmem2_6_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_6_ARLEN
        .m_axi_gmem2_6_ARSIZE   ( m_axi_gmem2_6_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_6_ARSIZE
        .m_axi_gmem2_6_ARBURST  ( m_axi_gmem2_6_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_6_ARBURST
        .m_axi_gmem2_6_ARLOCK   ( m_axi_gmem2_6_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_6_ARLOCK
        .m_axi_gmem2_6_ARREGION ( m_axi_gmem2_6_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_6_ARREGION
        .m_axi_gmem2_6_ARCACHE  ( m_axi_gmem2_6_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_6_ARCACHE
        .m_axi_gmem2_6_ARPROT   ( m_axi_gmem2_6_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_6_ARPROT
        .m_axi_gmem2_6_ARQOS    ( m_axi_gmem2_6_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_6_ARQOS
        .m_axi_gmem2_6_ARVALID  ( m_axi_gmem2_6_ARVALID  ) , // output wire m_axi_gmem2_6_ARVALID
        .m_axi_gmem2_6_ARREADY  ( m_axi_gmem2_6_ARREADY  ) , // input wire m_axi_gmem2_6_ARREADY
        .m_axi_gmem2_6_RDATA    ( m_axi_gmem2_6_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_6_RDATA
        .m_axi_gmem2_6_RRESP    ( m_axi_gmem2_6_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_6_RRESP
        .m_axi_gmem2_6_RLAST    ( m_axi_gmem2_6_RLAST    ) , // input wire m_axi_gmem2_6_RLAST
        .m_axi_gmem2_6_RVALID   ( m_axi_gmem2_6_RVALID   ) , // input wire m_axi_gmem2_6_RVALID
        .m_axi_gmem2_6_RREADY   ( m_axi_gmem2_6_RREADY   ) , // output wire m_axi_gmem2_6_RREADY
        .m_axi_gmem2_7_AWADDR   ( m_axi_gmem2_7_AWADDR   ) , // output wire [63 : 0] m_axi_gmem2_7_AWADDR
        .m_axi_gmem2_7_AWLEN    ( m_axi_gmem2_7_AWLEN    ) , // output wire [7 : 0] m_axi_gmem2_7_AWLEN
        .m_axi_gmem2_7_AWSIZE   ( m_axi_gmem2_7_AWSIZE   ) , // output wire [2 : 0] m_axi_gmem2_7_AWSIZE
        .m_axi_gmem2_7_AWBURST  ( m_axi_gmem2_7_AWBURST  ) , // output wire [1 : 0] m_axi_gmem2_7_AWBURST
        .m_axi_gmem2_7_AWLOCK   ( m_axi_gmem2_7_AWLOCK   ) , // output wire [1 : 0] m_axi_gmem2_7_AWLOCK
        .m_axi_gmem2_7_AWREGION ( m_axi_gmem2_7_AWREGION ) , // output wire [3 : 0] m_axi_gmem2_7_AWREGION
        .m_axi_gmem2_7_AWCACHE  ( m_axi_gmem2_7_AWCACHE  ) , // output wire [3 : 0] m_axi_gmem2_7_AWCACHE
        .m_axi_gmem2_7_AWPROT   ( m_axi_gmem2_7_AWPROT   ) , // output wire [2 : 0] m_axi_gmem2_7_AWPROT
        .m_axi_gmem2_7_AWQOS    ( m_axi_gmem2_7_AWQOS    ) , // output wire [3 : 0] m_axi_gmem2_7_AWQOS
        .m_axi_gmem2_7_AWVALID  ( m_axi_gmem2_7_AWVALID  ) , // output wire m_axi_gmem2_7_AWVALID
        .m_axi_gmem2_7_AWREADY  ( m_axi_gmem2_7_AWREADY  ) , // input wire m_axi_gmem2_7_AWREADY
        .m_axi_gmem2_7_WDATA    ( m_axi_gmem2_7_WDATA    ) , // output wire [63 : 0] m_axi_gmem2_7_WDATA
        .m_axi_gmem2_7_WSTRB    ( m_axi_gmem2_7_WSTRB    ) , // output wire [7 : 0] m_axi_gmem2_7_WSTRB
        .m_axi_gmem2_7_WLAST    ( m_axi_gmem2_7_WLAST    ) , // output wire m_axi_gmem2_7_WLAST
        .m_axi_gmem2_7_WVALID   ( m_axi_gmem2_7_WVALID   ) , // output wire m_axi_gmem2_7_WVALID
        .m_axi_gmem2_7_WREADY   ( m_axi_gmem2_7_WREADY   ) , // input wire m_axi_gmem2_7_WREADY
        .m_axi_gmem2_7_BRESP    ( m_axi_gmem2_7_BRESP    ) , // input wire [1 : 0] m_axi_gmem2_7_BRESP
        .m_axi_gmem2_7_BVALID   ( m_axi_gmem2_7_BVALID   ) , // input wire m_axi_gmem2_7_BVALID
        .m_axi_gmem2_7_BREADY   ( m_axi_gmem2_7_BREADY   ) , // output wire m_axi_gmem2_7_BREADY
        .m_axi_gmem2_7_ARADDR   ( m_axi_gmem2_7_ARADDR   ) , // output wire [63 : 0] m_axi_gmem2_7_ARADDR
        .m_axi_gmem2_7_ARLEN    ( m_axi_gmem2_7_ARLEN    ) , // output wire [7 : 0] m_axi_gmem2_7_ARLEN
        .m_axi_gmem2_7_ARSIZE   ( m_axi_gmem2_7_ARSIZE   ) , // output wire [2 : 0] m_axi_gmem2_7_ARSIZE
        .m_axi_gmem2_7_ARBURST  ( m_axi_gmem2_7_ARBURST  ) , // output wire [1 : 0] m_axi_gmem2_7_ARBURST
        .m_axi_gmem2_7_ARLOCK   ( m_axi_gmem2_7_ARLOCK   ) , // output wire [1 : 0] m_axi_gmem2_7_ARLOCK
        .m_axi_gmem2_7_ARREGION ( m_axi_gmem2_7_ARREGION ) , // output wire [3 : 0] m_axi_gmem2_7_ARREGION
        .m_axi_gmem2_7_ARCACHE  ( m_axi_gmem2_7_ARCACHE  ) , // output wire [3 : 0] m_axi_gmem2_7_ARCACHE
        .m_axi_gmem2_7_ARPROT   ( m_axi_gmem2_7_ARPROT   ) , // output wire [2 : 0] m_axi_gmem2_7_ARPROT
        .m_axi_gmem2_7_ARQOS    ( m_axi_gmem2_7_ARQOS    ) , // output wire [3 : 0] m_axi_gmem2_7_ARQOS
        .m_axi_gmem2_7_ARVALID  ( m_axi_gmem2_7_ARVALID  ) , // output wire m_axi_gmem2_7_ARVALID
        .m_axi_gmem2_7_ARREADY  ( m_axi_gmem2_7_ARREADY  ) , // input wire m_axi_gmem2_7_ARREADY
        .m_axi_gmem2_7_RDATA    ( m_axi_gmem2_7_RDATA    ) , // input wire [63 : 0] m_axi_gmem2_7_RDATA
        .m_axi_gmem2_7_RRESP    ( m_axi_gmem2_7_RRESP    ) , // input wire [1 : 0] m_axi_gmem2_7_RRESP
        .m_axi_gmem2_7_RLAST    ( m_axi_gmem2_7_RLAST    ) , // input wire m_axi_gmem2_7_RLAST
        .m_axi_gmem2_7_RVALID   ( m_axi_gmem2_7_RVALID   ) , // input wire m_axi_gmem2_7_RVALID
        .m_axi_gmem2_7_RREADY   ( m_axi_gmem2_7_RREADY   )   // output wire m_axi_gmem2_7_RREADY
    );

endmodule
